77330000 00090000 comctl32.dll
0fda0000 00030000 sccbase.dll
0fdd0000 00050000 slbcsp.dll
0fe20000 00180000 gpkcsp.dll
0ff80000 00020000 vdmredir.dll
0ff80000 000b0000 ntvdm.exe
0ffa0000 00010000 vcdex.dll
0ffa0000 00030000 dssenh.dll
0ffb0000 00050000 wow32.dll
0ffd0000 00030000 rsaenh.dll
47c80000 00010000 zextens.dll
47c90000 00010000 winclip.dll
47cb0000 00020000 ulkd.dll
47cd0000 00040000 traceprt.dll
47d10000 00020000 timerw32.dll
47d30000 00010000 statw32.dll
47d40000 00010000 secedt.dll
47d50000 00020000 sdbapiu.dll
47d70000 00020000 sdbapi.dll
47d90000 00020000 rwwin32.dll
47db0000 00010000 rwwin16.dll
47dc0000 00020000 rwres32.dll
47de0000 00020000 rwmac.dll
47e00000 00010000 rwinf.dll
47e20000 00010000 rcdata1.dll
47e30000 00010000 pptpkdx.dll
47e40000 00030000 ndrexts.dll
47e70000 00010000 nclipps.dll
47e80000 00040000 msiauto.dll
47ec0000 00010000 mepparty.dll
47ed0000 00020000 lsaexts.dll
47ef0000 00010000 irdakdx.dll
47f00000 00010000 iodll.dll
47f10000 00010000 dtext.dll
47f20000 00010000 depends.dll
47f30000 00010000 cxxflt.dll
47f40000 00010000 certexts.dll
47f50000 00010000 autosock.dll
47f60000 00020000 apidll.dll
47fb0000 00050000 adsiedit.dll
4be40000 00010000 wst.dll
4be90000 00010000 ulcase.dll
4bea0000 00010000 tglcase.dll
4beb0000 00010000 setupexts.dll
4bec0000 00010000 redbook.dll
4bed0000 00010000 pmatch.dll
4bee0000 00040000 msjvc.dll
4bf20000 00010000 mshelp.dll
4bf30000 00010000 mhelp.dll
4bf40000 00010000 justify.dll
4bf50000 00020000 jps.dll
4bf80000 00030000 iviewers.dll
4bfb0000 00030000 hwdll.dll
4bfe0000 00010000 filter.dll
4bff0000 00010000 dflayout.dll
4fae0000 00010000 shlexts.dll
4fb00000 00070000 msvcrtd.dll
4fb70000 00020000 msvcr40d.dll
4fb90000 00020000 msvcirtd.dll
4fbb0000 000d0000 mfco42ud.dll
4fc80000 000d0000 mfco42d.dll
4fd50000 00010000 mfcn42ud.dll
4fd60000 00010000 mfcn42d.dll
4fd70000 00050000 mfcd42ud.dll
4fdc0000 00050000 mfcd42d.dll
4fe10000 000f0000 mfc42ud.dll
4ff00000 000f0000 mfc42d.dll
4fff0000 00010000 conexts.dll
58170000 00040000 unimdm.tsp
581b0000 00020000 remotesp.tsp
581d0000 00010000 ndptsp.tsp
581f0000 00010000 kmddsp.tsp
58200000 00010000 ipconf.tsp
58210000 00010000 hidphone.tsp
58220000 00050000 h323.tsp
58270000 00070000 wmvds32.ax
582e0000 00070000 wmv8ds32.ax
58350000 00010000 wiasf.ax
58360000 00010000 vbisurf.ax
58370000 00010000 psisrndr.ax
58380000 00020000 phdsext.ax
583a0000 00020000 msscds32.ax
583c0000 00010000 msdvbnp.ax
583d0000 00040000 msadds32.ax
58410000 00070000 mpg4ds32.ax
58480000 00030000 mpg2splt.ax
584b0000 00010000 ksxbar.ax
584c0000 00020000 kswdmcap.ax
584e0000 00010000 kstvtune.ax
58500000 00020000 ksproxy.ax
58530000 00030000 ivfsrc.ax
58560000 000e0000 ir41_32.ax
58640000 00010000 ipsink.ax
58650000 00040000 iac25_32.ax
58690000 00010000 g711codc.ax
586a0000 00010000 dshowext.ax
586b0000 00020000 camext30.ax
586e0000 00040000 camext20.ax
58720000 00020000 camexo20.ax
58740000 00010000 bdaplgin.ax
58750000 00010000 agcgauge.ax
58760000 00020000 acelpdec.ax
58780000 00010000 tssoft32.acm
58790000 00020000 sl_anet.acm
587b0000 00010000 msgsm32.acm
587c0000 00020000 msg723.acm
587e0000 00010000 msg711.acm
587f0000 00050000 msaud32.acm
58840000 00090000 l3codeca.acm
588d0000 00010000 imaadp32.acm
588e0000 00020000 wshom.ocx
58900000 00030000 wmp.ocx
58940000 00020000 wmidx.ocx
58960000 00020000 tdc.ocx
58980000 00040000 sysmon.ocx
589c0000 00070000 swflash.ocx
58a30000 00020000 proctexe.ocx
58a50000 00020000 msscript.ocx
58a70000 00020000 logui.ocx
58a90000 00020000 ieinfo5.ocx
58ab0000 00020000 dmview.ocx
58ad0000 00020000 dhtmled.ocx
58b00000 00030000 daxctle.ocx
58b30000 00020000 cnfgprts.ocx
58b50000 00050000 certwiz.ocx
58ba0000 00020000 certmap.ocx
58bc0000 00020000 asctrls.ocx
58be0000 00020000 timedate.cpl
58c00000 00010000 telephon.cpl
58c10000 00050000 sysdm.cpl
58c60000 00030000 sapi.cpl
58c90000 00030000 powercfg.cpl
58cc0000 00010000 nwc.cpl
58cd0000 00050000 nusrmgr.cpl
58d40000 00010000 ncpa.cpl
58d50000 000a0000 mmsys.cpl
58df0000 00040000 main.cpl
58e30000 00020000 liccpa.cpl
58e50000 00010000 keymgr.cpl
58e60000 00020000 joy.cpl
58e80000 00010000 irprops.cpl
58ea0000 00030000 intl.cpl
58ed0000 00050000 inetcpl.cpl
58f30000 00030000 hdwwiz.cpl
58f60000 00030000 desk.cpl
58f90000 00020000 access.cpl
58fb0000 00050000 msh263.drv
59000000 00030000 msh261.drv
59030000 00010000 xxpclru1.dll
59040000 00030000 xuim750.dll
59070000 00010000 xrxwbtmp.dll
59080000 00010000 xrxscnui.dll
59090000 00040000 xrxnui.dll
590d0000 00010000 xrxnpcl.dll
590e0000 00030000 xrpr6res.dll
59110000 00010000 xrpclres.dll
59120000 00010000 xrenm760.dll
59130000 00010000 xrenm750.dll
59140000 00010000 xpclres1.dll
59150000 00010000 xolehlp.dll
59160000 00010000 wzcdlg.dll
59180000 00030000 wuv3is.dll
591b0000 00010000 wupdinfo.dll
591c0000 00010000 wstdecod.dll
591d0000 00010000 wshsv.dll
591e0000 00010000 wshrm.dll
591f0000 00010000 wshirda.dll
59200000 00010000 wship6.dll
59210000 00010000 wshcon.dll
59220000 00010000 wshclus.dll
59230000 00010000 wshatm.dll
59240000 00090000 wsecedit.dll
592d0000 00010000 wp9res.dll
592e0000 00010000 wp24res.dll
592f0000 00010000 wowfaxui.dll
59300000 00010000 wowfax.dll
59310000 000d0000 wmvdmoe.dll
593e0000 00070000 wmvdmod.dll
59450000 00070000 wmv8dmod.dll
594d0000 00050000 wmstream.dll
59530000 00020000 wmsocm.dll
59550000 00020000 wmsdmoe.dll
59570000 00020000 wmsdmod.dll
59590000 00080000 wmpvis.dll
59620000 00160000 wmpui.dll
59780000 00020000 wmpshell.dll
597a0000 001f0000 wmploc.dll
59990000 00140000 wmpcore.dll
59ad0000 00040000 wmpcd.dll
59b20000 00040000 wmnetmgr.dll
59b60000 00030000 wmmutil.dll
59b90000 00050000 wmmres.dll
59bf0000 00060000 wmmfilt.dll
59c50000 00020000 wmitimep.dll
59c70000 00020000 wmisvc.dll
59c90000 00010000 wmiscmgr.dll
59cb0000 00010000 wmipsess.dll
59cc0000 00070000 wmiprvsd.dll
59d30000 00010000 wmiprop.dll
59d40000 00020000 wmipjobj.dll
59d60000 00020000 wmipiprt.dll
59d80000 00020000 wmipicmp.dll
59da0000 00030000 wmipdskq.dll
59dd0000 00010000 wmipdfs.dll
59de0000 00030000 wmipcima.dll
59e10000 00030000 wmidcprv.dll
59e40000 00020000 wmicookr.dll
59e60000 00020000 wmiaprpl.dll
59e80000 00010000 wmiapres.dll
59e90000 00010000 wmi2xml.dll
59ea0000 00010000 wmerrsve.dll
59ec0000 00010000 wmerrenu.dll
59ee0000 00010000 wmdmps.dll
59ef0000 00010000 wmdmlog.dll
59f00000 00050000 wmasf.dll
59f50000 00080000 wmadmoe.dll
59fd0000 00040000 wmadmod.dll
5a010000 00020000 wlbsprov.dll
5a030000 00010000 wlbsctrl.dll
5a040000 00010000 wisc10.dll
5a050000 00010000 winstrm.dll
5a060000 000a0000 winssnap.dll
5a100000 00010000 winsrpc.dll
5a110000 00050000 winsmon.dll
5a160000 00010000 winsmib.dll
5a170000 00020000 winsevnt.dll
5a190000 00010000 winsctrs.dll
5a270000 00020000 wsdueng.dll
5a290000 00010000 wsdu.dll
5a2b0000 00010000 vidupgrd.dll
5a2c0000 00010000 tscomp.dll
5a330000 00010000 tjupg.dll
5a350000 00010000 spxupgrd.dll
5a360000 00020000 eqnupgrd.dll
5a380000 00010000 dgrpupg.dll
5a390000 00010000 digpriup.dll
5a3a0000 00020000 digiupg.dll
5a3c0000 00010000 dgupgrd.dll
5a3d0000 00010000 ntdsupg.dll
5a3e0000 00020000 netupgrd.dll
5a410000 00010000 msmqcomp.dll
5a420000 00010000 snadlcug.dll
5a430000 00010000 ntsnaupg.dll
5a440000 00010000 ibmmgug.dll
5a450000 00010000 mdmshrup.dll
5a460000 00010000 inpupgrd.dll
5a470000 00010000 ftcomp.dll
5a480000 00010000 fsfilter.dll
5a490000 00010000 cluscomp.dll
5a4c0000 00010000 boscomp.dll
5a4d0000 00010000 apmupgrd.dll
5a4e0000 000d0000 winntbbu.dll
5a680000 00190000 winnt32u.dll
5a810000 00120000 winnt32a.dll
5a950000 00020000 hwdb.dll
5a990000 00010000 winmgmtr.dll
5a9a0000 00030000 wiavusd.dll
5a9d0000 00020000 wiavideo.dll
5a9f0000 00090000 wiashext.dll
5aa80000 00020000 wiascr.dll
5aaa0000 00020000 wiamsmud.dll
5aac0000 00020000 wiafbdrv.dll
5aae0000 00020000 wiadss.dll
5ab10000 00070000 wiadefui.dll
5ab90000 00030000 webvw.dll
5abc0000 00010000 webhits.dll
5abd0000 00020000 webclnt.dll
5abf0000 00020000 wbemupgd.dll
5ac10000 00010000 wbemperf.dll
5ac20000 00030000 wbemdisp.dll
5ac50000 00030000 wbemcntl.dll
5ac90000 00010000 wbemads.dll
5aca0000 00040000 wavemsp.dll
5ace0000 00010000 wamregps.dll
5acf0000 00010000 wamreg51.dll
5ad10000 00010000 wamreg.dll
5ad20000 00010000 wamps51.dll
5ad30000 00010000 wamps.dll
5ad40000 00020000 wam51.dll
5ad60000 00010000 wam.dll
5ad70000 00020000 wabimp.dll
5ad90000 00010000 wabfind.dll
5ada0000 00040000 wab32res.dll
5adf0000 00080000 wab32.dll
5ae70000 00080000 w95upgnt.dll
5aef0000 00010000 w95inf32.dll
5af00000 00010000 w3tp.dll
5af10000 00060000 w3svc.dll
5af70000 00010000 w3svapi.dll
5af80000 00010000 w3ssl.dll
5af90000 00010000 w3scfg.dll
5afa0000 00010000 w3isapi.dll
5afb0000 00020000 w3ext.dll
5afd0000 00010000 w3dt.dll
5afe0000 00010000 w3ctrs51.dll
5aff0000 00010000 w3ctrs.dll
5b000000 00010000 w3ctrlps.dll
5b010000 00050000 w3core.dll
5b060000 00010000 w3comlog.dll
5b070000 00010000 w3cache.dll
5b080000 00010000 vwipxspx.dll
5b090000 00020000 vssui.dll
5b0b0000 00010000 vss_ps.dll
5b0c0000 00010000 vmmreg32.dll
5b0d0000 00010000 vjoy.dll
5b0e0000 00030000 viewprov.dll
5b110000 000d0000 vgx.dll
5b1e0000 00010000 vfwwdm32.dll
5b200000 00050000 verifier.dll
5b250000 00010000 vdmdbg.dll
5b260000 00010000 vbssv.dll
5b270000 00040000 uxtheme.dll
5b2b0000 00010000 utildll.dll
5b2c0000 00010000 usrvpa.dll
5b2d0000 00010000 usrvoica.dll
5b2e0000 00010000 usrv80a.dll
5b2f0000 00040000 usrv42a.dll
5b330000 00010000 usrsvpia.dll
5b340000 00010000 usrsdpia.dll
5b350000 00020000 usrrtosa.dll
5b370000 00010000 usrlbva.dll
5b380000 00020000 usrfaxa.dll
5b3a0000 00060000 usrdtea.dll
5b400000 00020000 usrdpa.dll
5b420000 00020000 usrcoina.dll
5b440000 00010000 usrcntra.dll
5b460000 00020000 usbui.dll
5b480000 00040000 upnpui.dll
5b4c0000 00030000 upnphost.dll
5b4f0000 00030000 updprov.dll
5b520000 00050000 untfs.dll
5b570000 00020000 unimdmat.dll
5b590000 00010000 uniansi.dll
5b5a0000 00010000 umdmxfrm.dll
5b5b0000 00020000 umaxud32.dll
5b5d0000 00010000 umaxu40.dll
5b5e0000 00010000 umaxu22.dll
5b5f0000 00030000 umaxu12.dll
5b620000 00020000 umaxscan.dll
5b640000 00020000 umaxp60.dll
5b660000 00010000 umaxcam.dll
5b680000 00010000 umandlg.dll
5b690000 00050000 um54scan.dll
5b6e0000 00050000 um34scan.dll
5b730000 00020000 uihelper.dll
5b750000 00020000 ufat.dll
5b770000 00010000 udhisapi.dll
5b780000 00010000 ty2x4res.dll
5b790000 00020000 ty2x3res.dll
5b7b0000 00020000 txflog.dll
5b7d0000 00010000 twain_32.dll
5b7f0000 00010000 ttyui.dll
5b800000 00010000 ttyres.dll
5b810000 00010000 tty.dll
5b820000 00010000 tsuserex.dll
5b830000 00010000 tssdjet.dll
5b840000 00020000 tsoc.dll
5b860000 00050000 tshoot.dll
5b8b0000 00010000 tsec.dll
5b8c0000 00020000 tscfgwmi.dll
5b8e0000 00050000 tscc.dll
5b930000 00010000 tsappcmp.dll
5b950000 00010000 trustmon.dll
5b960000 00020000 trnsprov.dll
5b980000 00010000 trksvr.dll
5b9a0000 00030000 triedit.dll
5b9d0000 00090000 tridxp.dll
5ba60000 00010000 trialoc.dll
5ba70000 00010000 tp4res.dll
5ba80000 00010000 tp4.dll
5ba90000 00010000 tools.dll
5baa0000 00020000 tmplprov.dll
5bac0000 00010000 tlyp6res.dll
5bad0000 00010000 tly5cres.dll
5bae0000 00010000 tly3res.dll
5bb00000 00010000 tls236.dll
5bb10000 00010000 tlntsvrp.dll
5bb20000 00010000 ti850res.dll
5bb30000 00080000 themeui.dll
5bbb0000 00030000 thawbrkr.dll
5bbf0000 00060000 termmgr.dll
5bc50000 00010000 tcpmonui.dll
5bc60000 00010000 tcdata.dll
5bc70000 00020000 tapiui.dll
5bc90000 00050000 tapisnap.dll
5bce0000 00010000 tapiperf.dll
5bcf0000 000d0000 tapi3.dll
5bdc0000 000f0000 t5000uni.dll
5beb0000 00010000 t5000ui.dll
5bed0000 00010000 t5000.dll
5bee0000 00010000 t3016.dll
5bef0000 000f0000 syssetup.dll
5bfe0000 00030000 sysmod_a.dll
5c010000 00030000 sysmod.dll
5c040000 00010000 sysinv.dll
5c050000 00010000 synceng.dll
5c070000 00020000 sxports.dll
5c0c0000 00010000 swpidflt.dll
5c0d0000 00010000 swpdflt2.dll
5c0e0000 00010000 sw_wheel.dll
5c100000 00010000 sw_effct.dll
5c110000 00010000 svcpack.dll
5c120000 00010000 svcext51.dll
5c130000 00010000 svcext.dll
5c150000 00010000 strmfilt.dll
5c160000 00040000 strmdll.dll
5c1b0000 00010000 streamci.dll
5c1c0000 00010000 str9eres.dll
5c1d0000 00020000 str24res.dll
5c1f0000 00020000 storprop.dll
5c210000 00030000 stlnprop.dll
5c240000 00010000 stlncoin.dll
5c250000 00010000 stjtres.dll
5c260000 00030000 sti_ci.dll
5c290000 00020000 stdprov.dll
5c2b0000 00020000 stclient.dll
5c2d0000 00010000 staxmem.dll
5c2e0000 00010000 status.dll
5c2f0000 00020000 star9res.dll
5c310000 00040000 st24eres.dll
5c360000 00010000 sstub.dll
5c370000 00010000 sspifilt.dll
5c380000 00010000 sslcfg.dll
5c390000 00010000 ssinc51.dll
5c3a0000 00010000 ssinc.dll
5c450000 00040000 swprv.dll
5c4e0000 00020000 srusd.dll
5c500000 00020000 srusbusd.dll
5c520000 00040000 srrstr.dll
5c560000 00020000 srclient.dll
5c580000 000d0000 srchui.dll
5c650000 00020000 srchctls.dll
5c670000 00040000 sqlxmlx.dll
5c6b0000 00030000 sqlunirl.dll
5c6e0000 00010000 spxupchk.dll
5c6f0000 00010000 spxcoins.dll
5c700000 000c0000 spttseng.dll
5c7c0000 00050000 sptip.dll
5c810000 00020000 sprio800.dll
5c830000 00020000 sprio600.dll
5c850000 00020000 spnike.dll
5c870000 00020000 spdports.dll
5c890000 00010000 spcplui.dll
5c8b0000 00020000 spcommon.dll
5c8d0000 00020000 sonypi.dll
5c900000 00020000 sonync.dll
5c930000 00030000 softkbd.dll
5c960000 00010000 snmpthrd.dll
5c970000 00010000 snmpstup.dll
5c980000 00030000 snmpsnap.dll
5c9c0000 00030000 snmpsmir.dll
5ca00000 00010000 snmpmib.dll
5ca10000 00060000 snmpincl.dll
5ca70000 00040000 snmpcl.dll
5cac0000 00010000 sniffpol.dll
5cad0000 00050000 snapshot.dll
5cb20000 00010000 smtpcons.dll
5cb30000 00020000 sml8xres.dll
5cb60000 00010000 smimsgif.dll
5cb70000 00010000 smierrsy.dll
5cb80000 00010000 smierrsm.dll
5cb90000 00010000 smb6w.dll
5cba0000 00010000 smb3w.dll
5cbb0000 00010000 smb0w.dll
5cbc0000 00010000 sma3w.dll
5cbd0000 00010000 sma0w.dll
5cbe0000 00010000 sm9aw.dll
5cbf0000 00010000 sm93w.dll
5cc00000 00010000 sm92w.dll
5cc10000 00010000 sm91w.dll
5cc20000 00010000 sm90w.dll
5cc30000 00010000 sm8dw.dll
5cc40000 00010000 sm8cw.dll
5cc50000 00010000 sm8aw.dll
5cc60000 00010000 sm89w.dll
5cc70000 00010000 sm87w.dll
5cc80000 00010000 sm81w.dll
5cc90000 00010000 sm59w.dll
5cca0000 00010000 slbs.dll
5ccb0000 00010000 slbrccsp.dll
5ccc0000 00020000 slbiop.dll
5cce0000 00010000 slayerxp.dll
5ccf0000 00010000 skdll.dll
5cd00000 00010000 skcolres.dll
5cd10000 00040000 sisgrv.dll
5cd50000 00010000 sisbkup.dll
5cd60000 00010000 simptcp.dll
5cd70000 00010000 sigtab.dll
5cd80000 00220000 shvlres.dll
5cfa0000 00020000 shvl.dll
5cfc0000 00010000 shscrap.dll
5cfd0000 00030000 shmedia.dll
5d000000 00070000 shimgvw.dll
5d070000 00030000 shimeng.dll
5d0a0000 00020000 sfmwshat.dll
5d0c0000 00010000 sfmpsprt.dll
5d0d0000 00010000 sfmpsfnt.dll
5d0e0000 000a0000 sfmpsdib.dll
5d190000 00010000 sfmmsg.dll
5d1a0000 00010000 sfmmon.dll
5d1b0000 00010000 sfmctrs.dll
5d1c0000 00010000 sfmatmsg.dll
5d1d0000 00010000 sfmapi.dll
5d1e0000 00020000 setupqry.dll
5d200000 00070000 setupdll.dll
5d270000 00010000 serwvdrv.dll
5d280000 00010000 servdeps.dll
5d2a0000 00010000 serialui.dll
5d2b0000 00010000 senscfg.dll
5d2c0000 00010000 sendmail.dll
5d2e0000 00010000 sendcmsg.dll
5d2f0000 00010000 sek9res.dll
5d300000 00010000 sek24res.dll
5d310000 00030000 sdpblb.dll
5d340000 00010000 scrrnsv.dll
5d350000 00030000 scrobj.dll
5d380000 00010000 scriptpw.dll
5d390000 00010000 scripto.dll
5d3a0000 00030000 script_a.dll
5d3d0000 00040000 script.dll
5d410000 00010000 scredir.dll
5d420000 00010000 scosv.dll
5d430000 00010000 sclgntfy.dll
5d440000 00030000 schmmgmt.dll
5d470000 00030000 sceprov.dll
5d4a0000 00030000 sccsccp.dll
5d4d0000 00020000 scardssp.dll
5d500000 00020000 scarddlg.dll
5d520000 00090000 sblfx.dll
5d5b0000 000b0000 sapi.dll
5d660000 00010000 safrslv.dll
5d670000 00010000 safrdm.dll
5d680000 00010000 safrcdlg.dll
5d690000 00020000 rwia450.dll
5d6b0000 00020000 rwia430.dll
5d6d0000 00020000 rwia330.dll
5d6f0000 00020000 rwia001.dll
5d710000 00010000 rw450ext.dll
5d720000 00010000 rw430ext.dll
5d730000 00010000 rw330ext.dll
5d740000 00010000 rw001ext.dll
5d750000 000c0000 rvseres.dll
5d810000 00010000 rvse.dll
5d830000 00010000 rtrupg.dll
5d840000 00020000 rtrfiltr.dll
5d860000 00020000 rtm.dll
5d880000 00010000 rtipxmib.dll
5d890000 00090000 rtcdll.dll
5d920000 00010000 rsvpperf.dll
5d930000 00010000 rsvpmsg.dll
5d940000 00060000 rstask.dll
5d9a0000 00010000 rssubps.dll
5d9b0000 00080000 rssub.dll
5da30000 00010000 rsshell.dll
5da40000 00010000 rsservps.dll
5da50000 00020000 rsoptcom.dll
5da70000 00010000 rsmps.dll
5da80000 00050000 rsmover.dll
5dad0000 00010000 rsmgrstr.dll
5dae0000 00090000 rsjob.dll
5db70000 00030000 rsidb.dll
5dba0000 00010000 rshx32.dll
5dbb0000 00010000 rsfsaps.dll
5dbc0000 00080000 rsfsa.dll
5dc40000 00010000 rsengps.dll
5dc50000 00030000 rseng.dll
5dc80000 00010000 rsconn.dll
5dc90000 00070000 rscommon.dll
5dd00000 00020000 rscli.dll
5dd30000 000e0000 rsadmin.dll
5de10000 00010000 rrasprxy.dll
5de20000 00010000 rpcref.dll
5de30000 00010000 rpcproxy.dll
5de40000 00010000 rpcns4.dll
5de50000 00010000 routetab.dll
5de60000 00010000 ripagnt.dll
5de70000 00010000 rigpsnap.dll
5de80000 00030000 ricohres.dll
5deb0000 00010000 riafui2.dll
5dec0000 00010000 riafui1.dll
5ded0000 00030000 riafres.dll
5df00000 00020000 reslog32.dll
5df20000 00010000 replprov.dll
5df30000 00020000 rend.dll
5df50000 00020000 remotepg.dll
5df70000 00070000 regwizc.dll
5dfe0000 00010000 rdpsnd.dll
5dff0000 00010000 rdpcfgex.dll
5e000000 00030000 rdchost.dll
5e030000 00020000 rcbdyctl.dll
5e050000 00030000 rasuser.dll
5e080000 00010000 rassfm.dll
5e090000 00010000 rasser.dll
5e0a0000 00010000 rasrad.dll
5e0b0000 00010000 rasmxs.dll
5e0c0000 00030000 rasmontr.dll
5e0f0000 00050000 rasdlg4.dll
5e140000 00010000 rasctrs.dll
5e150000 00010000 rasaudio.dll
5e160000 00010000 racpldlg.dll
5e170000 00010000 qvusd.dll
5e180000 00050000 msnsspc.dll
5e1d0000 00050000 wscsvc.dll
5e220000 000b0000 OPEN
5e2d0000 00010000 qosname.dll
5e2e0000 00010000 qmgrprxy.dll
5e2f0000 00050000 qmgr.dll
5e350000 000c0000 qedwipes.dll
5e410000 00080000 qedit.dll
5e4a0000 00060000 qdvd.dll
5e500000 00050000 qdv.dll
5e550000 00030000 qasf.dll
5e580000 00010000 pwsdata.dll
5e590000 00010000 pwdssp.dll
5e5a0000 00030000 ptpusd.dll
5e5d0000 00010000 ptpusb.dll
5e5e0000 00010000 pstorec.dll
5e5f0000 00010000 psnppagn.dll
5e600000 00010000 psisload.dll
5e610000 00070000 psisdecd.dll
5e680000 00080000 pscript5.dll
5e700000 00010000 pschdprf.dll
5e710000 00030000 ps5ui.dll
5e740000 00040000 provthrd.dll
5e780000 00080000 proccon.dll
5e800000 00010000 prflbmsg.dll
5e810000 00020000 policman.dll
5e830000 00010000 pngfilt.dll
5e840000 00200000 pmxviceo.dll
5ea40000 00010000 pmxmcro.dll
5ea50000 000d0000 pmxgl.dll
5eb20000 00010000 plustab.dll
5eb30000 00010000 plotui.dll
5eb50000 00010000 plotter.dll
5eb60000 00010000 pifmgr.dll
5eb80000 00010000 pid.dll
5eb90000 00030000 phvfwext.dll
5ebc0000 00030000 photowiz.dll
5ebf0000 00010000 philcam1.dll
5ec00000 00010000 permchk.dll
5ec60000 00010000 perfts.dll
5ec70000 00010000 perfproc.dll
5ec80000 00010000 perfos.dll
5ec90000 00010000 perfnw.dll
5eca0000 00010000 perfnet.dll
5ecb0000 00010000 perfdisk.dll
5ecc0000 00010000 perfctrs.dll
5ecd0000 00030000 pclxl.dll
5ed00000 00010000 pcleures.dll
5ed20000 000b0000 pcl5ures.dll
5edd0000 00040000 pcl4res.dll
5ee20000 00020000 pchshell.dll
5ee40000 00010000 pbsvrmsg.dll
5ee50000 00010000 pbsmon.dll
5ee60000 00010000 pbserver.dll
5ee70000 00020000 pautoenr.dll
5ee90000 00010000 parser.dll
5eea0000 00030000 paqsp.dll
5eed0000 00010000 panmap.dll
5eee0000 00010000 pagecnt.dll
5eef0000 00010000 pa9w9x.dll
5ef00000 00010000 pa9res.dll
5ef20000 00010000 pa24w9x.dll
5ef30000 00020000 pa24res.dll
5ef50000 000f0000 p5000uni.dll
5f040000 00010000 p5000ui.dll
5f050000 00010000 p5000.dll
5f060000 00010000 ovui2rc.dll
5f070000 00010000 ovui2.dll
5f080000 00010000 ovcomc.dll
5f090000 00020000 ovcodec2.dll
5f0c0000 00020000 osuninst.dll
5f0e0000 00020000 ospfmib.dll
5f100000 00010000 ospfagnt.dll
5f110000 00030000 ospf.dll
5f140000 00070000 optrares.dll
5f1b0000 00070000 opteures.dll
5f220000 000d0000 opengl32.dll
5f2f0000 00020000 olepro32.dll
5f310000 00020000 oleprn.dll
5f330000 00010000 oleaccrc.dll
5f340000 00010000 old9res.dll
5f350000 00010000 old24res.dll
5f360000 00010000 ol9res.dll
5f370000 00010000 ol24res.dll
5f380000 00010000 oksidm9.dll
5f390000 00030000 okml9res.dll
5f3c0000 00020000 okm24res.dll
5f3e0000 00030000 okipage.dll
5f410000 00010000 oki9res.dll
5f420000 00010000 oki24res.dll
5f430000 00010000 okd24res.dll
5f450000 00020000 ok9ibres.dll
5f470000 00020000 offfilt.dll
5f490000 00010000 oemiglib.dll
5f4a0000 00020000 oeimport.dll
5f4c0000 00010000 odbcp32r.dll
5f4d0000 00020000 odbcconf.dll
5f500000 00020000 od9ibres.dll
5f520000 00010000 ocmsn.dll
5f530000 00020000 ocmanage.dll
5f550000 00010000 ocgen.dll
5f560000 00010000 oce.dll
5f570000 00020000 occache.dll
5f590000 00050000 objsel.dll
5f5e0000 00020000 nwwks.dll
5f600000 00030000 nwprovau.dll
5f630000 00010000 nwevent.dll
5f640000 00010000 nwcfg.dll
5f650000 00020000 nwapi32.dll
5f670000 00010000 nwapi16.dll
5f680000 00010000 ntvdmd.dll
5f690000 00010000 ntsdexts.dll
5f6a0000 00020000 ntprint.dll
5f6c0000 00020000 ntoc.dll
5f6e0000 00010000 ntmsevt.dll
5f6f0000 00010000 ntlanui2.dll
5f700000 00020000 ntfrsres.dll
5f720000 00010000 ntfrsprf.dll
5f730000 00010000 ntfrsapi.dll
5f750000 00040000 ntevt.dll
5f790000 00010000 ntdsperf.dll
5f7a0000 00060000 ntdsmsg.dll
5f800000 00010000 ntdsbmsg.dll
5f810000 00010000 nsepm.dll
5f820000 00010000 npwmsdrm.dll
5f830000 00010000 npptools.dll
5f850000 00060000 npdsplay.dll
5f8b0000 00030000 rsaenhs.dll
5f8e0000 00030000 nmwb.dll
5f910000 00010000 nmsupp.dll
5f920000 00010000 nmpppoe.dll
5f930000 00030000 nmoldwb.dll
5f960000 00010000 nmmkcert.dll
5f970000 00030000 nmft.dll
5f9a0000 00010000 nmevtmsg.dll
5f9b0000 00020000 nmapi.dll
5f9d0000 00020000 nlhtml.dll
5f9f0000 00030000 nlbmprov.dll
5fa20000 00010000 nextlink.dll
5fa40000 00040000 newdev.dll
5fa80000 000e0000 netplwiz.dll
5fb60000 00020000 netoc.dll
5fb80000 00030000 netid.dll
5fbb0000 00040000 neth.dll
5fc00000 00010000 ndisnpp.dll
5fc20000 00010000 nddenb32.dll
5fc30000 00010000 ncxpnt.dll
5fc40000 00010000 ncpsui.dll
5fc50000 00010000 ncpsres.dll
5fc60000 00020000 ncprov.dll
5fc80000 00010000 ncpclres.dll
5fc90000 00010000 ncobjapi.dll
5fca0000 00010000 nc24res.dll
5fcb0000 00020000 narrhook.dll
5fcd0000 000c0000 napmmc.dll
5fd90000 00010000 mxport.dll
5fda0000 00010000 mxicfg.dll
5fdb0000 00020000 mwci32.dll
5fdd0000 00010000 mty9res.dll
5fde0000 00030000 mty24res.dll
5fe10000 00010000 mtxlegih.dll
5fe20000 00010000 mtxex.dll
5fe30000 00010000 mtxdm.dll
5fe40000 00030000 mtpclres.dll
5fe70000 00010000 mtltres.dll
5fe80000 00010000 mtbjres.dll
5fe90000 00010000 mt90res.dll
5fea0000 00010000 mt735res.dll
5feb0000 00010000 msxmlr.dll
5fec0000 00010000 msxml3r.dll
5fed0000 00010000 msxml2r.dll
5fee0000 000b0000 msxml2.dll
5ff90000 00030000 mswmdm.dll
5ffc0000 00040000 mswebdvd.dll
5fff0000 00010000 kbd101.dll
5fff0000 00010000 kbd101a.dll
5fff0000 00010000 kbd101b.dll
5fff0000 00010000 kbd101c.dll
5fff0000 00010000 kbd103.dll
5fff0000 00010000 kbd106.dll
5fff0000 00010000 kbd106n.dll
5fff0000 00010000 kbdal.dll
5fff0000 00010000 kbdarme.dll
5fff0000 00010000 kbdarmw.dll
5fff0000 00010000 kbdax2.dll
5fff0000 00010000 kbdaze.dll
5fff0000 00010000 kbdazel.dll
5fff0000 00010000 kbdbe.dll
5fff0000 00010000 kbdbene.dll
5fff0000 00010000 kbdblr.dll
5fff0000 00010000 kbdbr.dll
5fff0000 00010000 kbdbu.dll
5fff0000 00010000 kbdca.dll
5fff0000 00010000 kbdcan.dll
5fff0000 00010000 kbdcr.dll
5fff0000 00010000 kbdcz.dll
5fff0000 00010000 kbdcz1.dll
5fff0000 00010000 kbdcz2.dll
5fff0000 00010000 kbdda.dll
5fff0000 00010000 kbddv.dll
5fff0000 00010000 kbdes.dll
5fff0000 00010000 kbdest.dll
5fff0000 00010000 kbdfc.dll
5fff0000 00010000 kbdfi.dll
5fff0000 00010000 kbdfo.dll
5fff0000 00010000 kbdfr.dll
5fff0000 00010000 kbdgae.dll
5fff0000 00010000 kbdgeo.dll
5fff0000 00010000 kbdgkl.dll
5fff0000 00010000 kbdgr.dll
5fff0000 00010000 kbdgr1.dll
5fff0000 00010000 kbdhe.dll
5fff0000 00010000 kbdhe220.dll
5fff0000 00010000 kbdhe319.dll
5fff0000 00010000 kbdhela2.dll
5fff0000 00010000 kbdhela3.dll
5fff0000 00010000 kbdhept.dll
5fff0000 00010000 kbdhu.dll
5fff0000 00010000 kbdhu1.dll
5fff0000 00010000 kbdibm02.dll
5fff0000 00010000 kbdic.dll
5fff0000 00010000 kbdir.dll
5fff0000 00010000 kbdit.dll
5fff0000 00010000 kbdit142.dll
5fff0000 00010000 kbdjpn.dll
5fff0000 00010000 kbdkaz.dll
5fff0000 00010000 kbdkor.dll
5fff0000 00010000 kbdla.dll
5fff0000 00010000 kbdlk41a.dll
5fff0000 00010000 kbdlk41j.dll
5fff0000 00010000 kbdlt.dll
5fff0000 00010000 kbdlt1.dll
5fff0000 00010000 kbdlv.dll
5fff0000 00010000 kbdlv1.dll
5fff0000 00010000 kbdmac.dll
5fff0000 00010000 kbdne.dll
5fff0000 00010000 kbdnec.dll
5fff0000 00010000 kbdnec95.dll
5fff0000 00010000 kbdnecat.dll
5fff0000 00010000 kbdnecnt.dll
5fff0000 00010000 kbdno.dll
5fff0000 00010000 kbdpl.dll
5fff0000 00010000 kbdpl1.dll
5fff0000 00010000 kbdpo.dll
5fff0000 00010000 kbdro.dll
5fff0000 00010000 kbdru.dll
5fff0000 00010000 kbdru1.dll
5fff0000 00010000 kbdsf.dll
5fff0000 00010000 kbdsg.dll
5fff0000 00010000 kbdsl.dll
5fff0000 00010000 kbdsl1.dll
5fff0000 00010000 kbdsp.dll
5fff0000 00010000 kbdsw.dll
5fff0000 00010000 kbdtat.dll
5fff0000 00010000 kbdtuf.dll
5fff0000 00010000 kbdtuq.dll
5fff0000 00010000 kbduk.dll
5fff0000 00010000 kbdur.dll
5fff0000 00010000 kbdus.dll
5fff0000 00010000 kbdusa.dll
5fff0000 00010000 kbdusl.dll
5fff0000 00010000 kbdusr.dll
5fff0000 00010000 kbdusx.dll
5fff0000 00010000 kbduzb.dll
5fff0000 00010000 kbdvntc.dll
5fff0000 00010000 kbdycc.dll
5fff0000 00010000 kbdycl.dll
60010000 00020000 msw3prt.dll
60030000 00100000 OPEN
60130000 00040000 msutb.dll
60170000 00040000 msuni11.dll
601b0000 00050000 mstvgs.dll
60200000 00060000 mstvca.dll
60260000 00030000 mstsmmc.dll
60290000 00020000 mstsmhst.dll
602b0000 00090000 OPEN
60340000 00080000 mstime.dll
603c0000 00010000 mst123.dll
603d0000 00010000 msswch.dll
603e0000 00010000 mssoapr.dll
603f0000 00040000 mssoap1.dll
60430000 00010000 mssip32.dll
60440000 00030000 msrating.dll
60470000 00020000 msratelc.dll
60490000 00010000 msr2cenu.dll
604a0000 00020000 msr2c.dll
604c0000 00010000 msppnxus.dll
604d0000 00040000 msppmgr.dll
60510000 00010000 msppmd5.dll
60520000 00010000 msppmalr.dll
60530000 00010000 mspplkrh.dll
60550000 00010000 msppcntr.dll
60560000 00010000 msppalrt.dll
60570000 00010000 msports.dll
60580000 00040000 mspmsp.dll
605c0000 00010000 mspatcha.dll
605d0000 00010000 msorc32r.dll
605e0000 00270000 msoeres.dll
60850000 00040000 msoeacct.dll
60890000 00130000 msoe.dll
609c0000 00010000 msobweb.dll
609d0000 00010000 msobshel.dll
609e0000 00090000 msobmain.dll
60a70000 00010000 msobjs.dll
60a80000 00010000 msobdl.dll
60a90000 00020000 msobcomm.dll
60ab0000 00030000 msmqocm.dll
60ae0000 00010000 mslwvtts.dll
60af0000 00010000 mslbui.dll
60b10000 00010000 msisip.dll
60b20000 00060000 msisam11.dll
60b80000 00050000 msiprov.dll
60bd0000 00060000 msinfo.dll
60c30000 000d0000 msimsg.dll
60d10000 00050000 msihnd.dll
60d70000 00040000 msieftp.dll
60db0000 00010000 msidntld.dll
60dc0000 00010000 msident.dll
60dd0000 00010000 mshtmler.dll
60df0000 00010000 msgrocm.dll
60e00000 00340000 msgr3en.dll
61140000 00020000 msencode.dll
61160000 00010000 msdxmlc.dll
61170000 00020000 msdvdopt.dll
61190000 00030000 msdtcuiu.dll
611c0000 000e0000 msdtctm.dll
612a0000 00020000 msdtcstp.dll
612c0000 00060000 msdtcprx.dll
61320000 00020000 msdtclog.dll
61340000 00010000 msdaurl.dll
61350000 00020000 msdatl3.dll
61370000 00010000 msdaprsr.dll
61380000 00010000 msdaorar.dll
61390000 00020000 msctfp.dll
613b0000 00010000 mscpx32r.dll
613c0000 00010000 msconf.dll
613e0000 00040000 msclus.dll
61420000 00040000 mscandui.dll
61460000 00020000 msaudite.dll
61480000 00020000 msaatext.dll
614a0000 00080000 mqutil.dll
61520000 00010000 mqupgrd.dll
61530000 00030000 mqtrig.dll
61560000 00010000 mqtgclus.dll
61570000 00080000 mqsnap.dll
615f0000 00020000 mqsec.dll
61610000 00020000 mqrtdep.dll
61640000 00030000 mqrt.dll
61670000 00010000 mqrperf.dll
61680000 000b0000 mqqm.dll
61730000 00010000 mqperf.dll
61740000 00040000 mqoa.dll
61780000 00040000 mqmigrat.dll
617c0000 00020000 mqlogmgr.dll
617e0000 00010000 mqise.dll
617f0000 00020000 mqgentr.dll
61810000 00010000 mqdssrv.dll
61820000 00010000 mqdscli.dll
61840000 00010000 mqdbodbc.dll
61850000 00020000 mqclus.dll
61870000 00010000 mqcertui.dll
61880000 00040000 mqads.dll
618c0000 00030000 mqad.dll
618f0000 00040000 mq1repl.dll
61930000 00100000 mprsnap.dll
61a30000 00020000 mprmsg.dll
61a50000 00010000 mprdim.dll
61a70000 00020000 mprddm.dll
61a90000 00060000 mpg4dmod.dll
61af0000 00040000 moricons.dll
61b30000 00020000 mofd.dll
61b60000 00010000 modex.dll
61b70000 00030000 modemui.dll
61ba0000 00040000 mobsync.dll
61be0000 00030000 mn350620.dll
61c10000 00030000 mmutilse.dll
61c40000 00010000 mmfutil.dll
61c50000 000a0000 mltres.dll
61cf0000 00010000 mll_qic.dll
61d00000 00010000 mll_mtf.dll
61d10000 00010000 mll_hp.dll
61d20000 00010000 miscanw.dll
61d30000 00040000 minqmsui.dll
61d70000 00010000 minqmsps.dll
61d80000 00030000 minolres.dll
61db0000 00030000 mindex.dll
61de0000 00010000 mimefilt.dll
61df0000 00020000 miglibnt.dll
61e10000 00040000 migism_a.dll
61e50000 00040000 migism.dll
61e90000 00020000 mga.dll
61eb0000 00010000 mfcsubs.dll
61ec0000 00010000 mfc42sve.dll
61ed0000 000f0000 mfc40u.dll
61fc0000 00010000 mfc40sve.dll
61fd0000 000f0000 mfc40.dll
620c0000 00060000 metal_ss.dll
62120000 00040000 metadata.dll
62160000 00020000 metada51.dll
62180000 00090000 memgrp.dll
62210000 00030000 mdwmdmsp.dll
62240000 00010000 mdsync.dll
62250000 00020000 mdminst.dll
62270000 00020000 mdhcp.dll
62290000 00010000 md5filt.dll
622a0000 00010000 mciwave.dll
622b0000 00010000 mciseq.dll
622c0000 00010000 mciqtz32.dll
622d0000 00010000 mciole32.dll
622e0000 00010000 mcicda.dll
62300000 00010000 mchgrcoi.dll
62310000 00010000 mcd32.dll
62320000 00010000 mcastmib.dll
62330000 00010000 mcast.dll
62340000 00020000 mapistub.dll
62370000 00010000 mag_hook.dll
62380000 00020000 m3092dc.dll
623a0000 00020000 m3091dc.dll
623c0000 00030000 lxsysui.dll
623f0000 00010000 lxsysres.dll
62400000 00010000 lxsysrdr.dll
62410000 00060000 lxsyicur.dll
62470000 00020000 lxsyfcic.dll
624a0000 000f0000 lxsdclr2.dll
62590000 001c0000 lxsdclr1.dll
62750000 00030000 lxrosui.dll
62780000 00010000 lxrosres.dll
62790000 00010000 lxrosrdr.dll
627a0000 00060000 lxroicur.dll
62800000 00020000 lxrofcic.dll
62830000 00030000 lxmdsui.dll
62860000 00010000 lxmdsres.dll
62870000 00010000 lxmdsrdr.dll
62880000 00060000 lxmdicur.dll
628e0000 00030000 lxmdfcic.dll
62910000 00030000 lxmasui.dll
62940000 00010000 lxmasres.dll
62950000 00010000 lxmasrdr.dll
62960000 00060000 lxmaicur.dll
629c0000 00020000 lxmafcic.dll
629f0000 00010000 lxinkres.dll
62a10000 00010000 lxfmpres.dll
62a20000 00030000 lxcasui.dll
62a50000 00010000 lxcasres.dll
62a60000 00010000 lxcasrdr.dll
62a70000 00060000 lxcaicur.dll
62ad0000 00030000 lxcafcic.dll
62b00000 00030000 lxaesui.dll
62b30000 00010000 lxaesres.dll
62b40000 00010000 lxaesrdr.dll
62b50000 00060000 lxaeicur.dll
62bb0000 00030000 lxaefcic.dll
62be0000 00030000 lxadsui.dll
62c10000 00010000 lxadsres.dll
62c20000 00010000 lxadsrdr.dll
62c30000 00060000 lxadicur.dll
62c90000 00030000 lxadfcic.dll
62cc0000 00030000 lxacsui.dll
62cf0000 00010000 lxacsres.dll
62d00000 00010000 lxacsrdr.dll
62d10000 00060000 lxacicur.dll
62d70000 00030000 lxacfcic.dll
62da0000 00030000 lxaasui.dll
62dd0000 00010000 lxaasres.dll
62de0000 00010000 lxaasrdr.dll
62df0000 00060000 lxaaicur.dll
62e50000 00030000 lxaafcic.dll
62e80000 00010000 lx238res.dll
62e90000 00040000 lrwizdll.dll
62ed0000 00010000 lprmonui.dll
62ee0000 00010000 lprmon.dll
62ef0000 00010000 lprhelp.dll
62f00000 00010000 lpk.dll
62f10000 00010000 lpdsvc.dll
62f20000 00010000 lonsint.dll
62f30000 00010000 logscrpt.dll
62f40000 00020000 loghours.dll
62f60000 00010000 log.dll
62f70000 00010000 localui.dll
62f80000 00060000 lmrt.dll
62ff0000 00030000 lmpclres.dll
63020000 00090000 lmoptra.dll
630b0000 00010000 lmmib2.dll
630c0000 00010000 lmikjres.dll
630d0000 00010000 llsrpc.dll
630f0000 00020000 licwmi.dll
63110000 00010000 licmgr10.dll
63120000 00010000 licenoc.dll
63130000 00060000 licdll.dll
63190000 00010000 lexutil.dll
631a0000 00010000 laprxy.dll
631b0000 00020000 langwrbk.dll
631d0000 00020000 voicesub.dll
631f0000 00110000 voicepad.dll
63300000 00020000 uniime.dll
63320000 00020000 tmigrate.dll
63340000 00030000 softkey.dll
63370000 00020000 pmigrate.dll
63390000 00020000 pintlcsd.dll
633b0000 00050000 pintlcsa.dll
63410000 00010000 padrs804.dll
63420000 00010000 padrs412.dll
63430000 00010000 padrs411.dll
63440000 00010000 padrs404.dll
63450000 00040000 multibox.dll
63490000 00020000 msir3jp.dll
634b0000 00020000 korwbrkr.dll
634d0000 00060000 imskf.dll
63530000 00080000 imskdic.dll
635b0000 00020000 imlang.dll
635d0000 00050000 imjputyc.dll
63620000 00020000 imjpdct.dll
63640000 000c0000 imjpcus.dll
63700000 00060000 imjpcic.dll
63760000 000d0000 imjp81k.dll
63830000 00020000 imepadsm.dll
63850000 00020000 imekrmbx.dll
63870000 00020000 imekrcic.dll
63890000 009b0000 hwxkor.dll
64240000 00ce0000 hwxjpn.dll
64f20000 009b0000 hwxcht.dll
658d0000 00010000 hanjadic.dll
658e0000 00010000 ftlx0411.dll
658f0000 00060000 cintime.dll
65950000 00060000 chtskf.dll
659b0000 00030000 chtskdic.dll
659e0000 00040000 chtmbx.dll
65a20000 000d0000 chtbrkr.dll
65b00000 001a0000 chsbrkr.dll
65ca0000 00020000 lamebtn.dll
65cc0000 00010000 kyrares.dll
65cd0000 00030000 kyores.dll
65d00000 00020000 kyofonts.dll
65d20000 00010000 krnlprov.dll
65d30000 00010000 kousd.dll
65d40000 00070000 kmres.dll
65db0000 00040000 keymgr.dll
65df0000 00010000 kerbprsr.dll
65e00000 00050000 kdsusd.dll
65e50000 00020000 kdsui.dll
65e80000 00030000 kdcsvc.dll
65eb0000 00010000 kbdurdu.dll
65ec0000 00010000 kbdth3.dll
65ed0000 00010000 kbdth2.dll
65ee0000 00010000 kbdth1.dll
65ef0000 00010000 kbdth0.dll
65f00000 00010000 kbdsyr2.dll
65f10000 00010000 kbdsyr1.dll
65f20000 00010000 kbdmon.dll
65f30000 00010000 kbdkyr.dll
65f40000 00010000 kbdintel.dll
65f50000 00010000 kbdintam.dll
65f60000 00010000 kbdinpun.dll
65f70000 00010000 kbdinmar.dll
65f80000 00010000 kbdinkan.dll
65f90000 00010000 kbdinhin.dll
65fa0000 00010000 kbdinguj.dll
65fb0000 00010000 kbdindev.dll
65fc0000 00010000 kbdheb.dll
65fd0000 00010000 kbdfa.dll
65fe0000 00010000 kbddiv2.dll
65ff0000 00010000 kbddiv1.dll
66000000 00010000 kbda3.dll
66010000 00010000 kbda2.dll
66020000 00010000 kbda1.dll
66030000 00010000 jupiw.dll
66040000 00010000 jssv.dll
66050000 00010000 jsproxy.dll
66060000 00020000 jp350res.dll
66090000 00010000 jobexec.dll
660b0000 00020000 jgsh400.dll
660d0000 00020000 jgsd400.dll
660f0000 00020000 jgpl400.dll
66110000 00010000 jgmd400.dll
66130000 00030000 jgdw400.dll
66160000 00010000 jgaw400.dll
66180000 000d0000 jet500.dll
66250000 000b0000 jet.dll
66300000 00010000 ixsso.dll
66320000 00010000 iwrps.dll
66330000 00030000 iuengine.dll
66360000 00020000 iuctl.dll
66380000 00030000 itss.dll
663b0000 00030000 itircl.dll
663e0000 00010000 isrdbg32.dll
663f0000 00010000 ismsmtp.dll
66410000 00010000 ismsink.dll
66420000 00010000 ismip.dll
66430000 00010000 ism.dll
66440000 00020000 isign32.dll
66460000 00010000 iscomlog.dll
66470000 00020000 isatq.dll
66490000 00010000 isapips.dll
664a0000 00020000 irmon.dll
664c0000 00010000 irclass.dll
664d0000 00090000 ir50_qc.dll
66560000 000b0000 ir41_qc.dll
66610000 00080000 ipxsnap.dll
66690000 00020000 ipxsap.dll
666b0000 00010000 ipxrtmgr.dll
666c0000 00010000 ipxrip.dll
666d0000 00020000 ipxpromn.dll
666f0000 00020000 ipxmontr.dll
66710000 00030000 ipv6mon.dll
66740000 000d0000 ipsnap.dll
66810000 00060000 ipsmsnap.dll
66870000 00060000 ipsecsnp.dll
668d0000 00030000 iprtrmgr.dll
66910000 00010000 iprtprio.dll
66920000 00010000 iprop.dll
66930000 00020000 iprip2.dll
66950000 00010000 iprip.dll
66960000 00060000 ippromon.dll
669c0000 00080000 ipnathlp.dll
66a40000 00030000 ipmontr.dll
66a70000 00010000 ipm.dll
66a80000 00010000 ipbootp.dll
66a90000 00010000 iologmsg.dll
66aa0000 00020000 io8ports.dll
66ac0000 00020000 inseng.dll
66ae0000 00020000 OPEN
66b00000 00030000 initpki.dll
66b30000 00080000 infosoft.dll
66bb0000 00010000 infoctrs.dll
66bc0000 00050000 infocomm.dll
66c10000 00010000 infoadmn.dll
66c20000 00010000 inetsloc.dll
66c30000 00010000 inetres.dll
66c40000 00010000 inetppui.dll
66c50000 00010000 inetmib1.dll
66c60000 000d0000 inetmgr.dll
66d30000 00020000 inetcplc.dll
66d50000 00050000 inetcfg.dll
66da0000 00030000 imsinsnt.dll
66dd0000 00010000 imirror.dll
66de0000 00010000 imgutil.dll
66df0000 00010000 imeshare.dll
66e00000 00020000 imadmui.dll
66e20000 00020000 ils.dll
66e40000 00030000 iiswmi.dll
66e70000 00020000 iisw3adm.dll
66e90000 00020000 iisutil.dll
66ec0000 00030000 iisui.dll
66f00000 00010000 iissuba.dll
66f10000 00020000 iisrtl.dll
66f40000 00010000 iisrstap.dll
66f50000 00010000 iismui.dll
66f60000 00020000 iismap.dll
66f80000 00020000 iislog51.dll
66fa0000 00020000 iislog.dll
66fc0000 00010000 iisfecnv.dll
66fd0000 00020000 iisext51.dll
66ff0000 00020000 iisext.dll
67010000 00010000 iiscrmap.dll
67020000 00010000 iisclus3.dll
67030000 00020000 iisclex4.dll
67050000 00020000 iisclex3.dll
67070000 00030000 iische51.dll
670a0000 001c0000 iiscfg.dll
67270000 00010000 iisadmin.dll
67280000 00080000 iis.dll
67300000 00030000 igmpv2.dll
67330000 00010000 igmpagnt.dll
67340000 00020000 ifsutil.dll
67360000 00030000 ifmon.dll
67390000 00020000 iesetup.dll
673b0000 00010000 iernonce.dll
673c0000 00040000 iepeers.dll
67400000 00050000 iedkcs32.dll
67450000 00040000 ieakui.dll
67490000 00040000 ieaksie.dll
674d0000 00020000 ieakeng.dll
67500000 00020000 idq.dll
67520000 00010000 icwutil.dll
67530000 00010000 icwres.dll
67550000 00010000 icwphbk.dll
67570000 00030000 icwhelp.dll
675a0000 00010000 icwdl.dll
675b0000 00020000 icwdial.dll
675d0000 00010000 icwconn.dll
675e0000 00010000 iconlib.dll
675f0000 00060000 iconf32.dll
67660000 00010000 icmui.dll
67680000 00040000 icm32.dll
676c0000 00010000 icfgnt5.dll
676d0000 00010000 icam5ext.dll
676e0000 00010000 icam5com.dll
676f0000 00020000 icam4ext.dll
67710000 00020000 icam4com.dll
67730000 00010000 icam3ext.dll
67740000 00010000 ibqwres.dll
67750000 00010000 ibps1res.dll
67760000 00010000 ibprores.dll
67770000 00010000 ibppdres.dll
67780000 00010000 ibp24res.dll
67790000 00010000 ibmsgnet.dll
677a0000 00010000 ibmptres.dll
677b0000 00010000 ib52res.dll
677c0000 00010000 ib239res.dll
677e0000 00010000 ib238res.dll
677f0000 00020000 iassvcs.dll
67810000 00040000 iassdo.dll
67860000 00020000 iassam.dll
67880000 00030000 iasrecst.dll
678b0000 00020000 iasrad.dll
678e0000 00010000 iaspolcy.dll
678f0000 00010000 iasperf.dll
67900000 00020000 iasnap.dll
67920000 00040000 iasmmc.dll
67970000 00010000 iashlpr.dll
67980000 00010000 iasads.dll
67990000 00010000 iasacct.dll
679a0000 00010000 ias.dll
679b0000 00080000 hypertrm.dll
67a30000 00010000 htui.dll
67a40000 00010000 httpodbc.dll
67a50000 00020000 httpod51.dll
67a70000 00010000 httpmib.dll
67a80000 00010000 httpmb51.dll
67a90000 00040000 httpext.dll
67ae0000 00010000 httpapi.dll
67af0000 00010000 htrn_jis.dll
67b00000 00010000 hsf_inst.dll
67b10000 00130000 hrtzres.dll
67c40000 00020000 hrtz.dll
67c60000 00010000 hr1w.dll
67c70000 00040000 hpwm5db1.dll
67cb0000 00050000 hpwm50al.dll
67d00000 00010000 hpvui50.dll
67d10000 00020000 hpvud50.dll
67d30000 00030000 hpvscp50.dll
67d70000 00280000 hpvimg50.dll
67ff0000 00040000 hpvdb820.dll
68030000 00030000 hpvdb720.dll
68060000 00080000 hpv880al.dll
680e0000 00050000 hpv850al.dll
68130000 00060000 hpv820al.dll
68190000 00050000 hpv800al.dll
681f0000 00060000 hpv700al.dll
68250000 00050000 hpv600al.dll
682a0000 00060000 hpv200al.dll
68300000 00010000 hptjres.dll
68310000 00010000 hpsjmcro.dll
68320000 00010000 hpqjres.dll
68330000 00010000 hppjres.dll
68340000 00060000 hpojwia.dll
683a0000 00010000 hpoemui.dll
683b0000 00010000 hpmcro32.dll
683c0000 00010000 hpgtmcro.dll
683d0000 00020000 hpgt53tk.dll
683f0000 00030000 hpgt53.dll
68420000 00010000 hpgt42tk.dll
68430000 00020000 hpgt42.dll
68450000 00150000 hpgt34tk.dll
685a0000 00020000 hpgt34.dll
685c0000 00140000 hpgt33tk.dll
68700000 00020000 hpgt33.dll
68720000 00030000 hpgt21tk.dll
68750000 00020000 hpgt21.dll
68770000 00010000 hpfui50.dll
68780000 00020000 hpfud50.dll
687a0000 001d0000 hpfimg50.dll
68970000 000e0000 hpf940al.dll
68a50000 00070000 hpf900al.dll
68ac0000 00080000 hpf880al.dll
68b40000 00030000 hpdjres.dll
68b70000 00030000 hpdigwia.dll
68ba0000 00010000 hpcstr.dll
68bb0000 00060000 hpclj5ui.dll
68c10000 00010000 hpcjrui.dll
68c20000 00010000 hpcjrrps.dll
68c30000 00010000 hpcjrr.dll
68c40000 00030000 hpcfont.dll
68c70000 00010000 hpccljui.dll
68c80000 00010000 hpcclj1.dll
68c90000 00010000 hpcclj.dll
68ca0000 00010000 hpcabout.dll
68cb0000 00020000 hpc4500u.dll
68ce0000 00030000 hotplug.dll
68d10000 00010000 hostmib.dll
68d20000 00060000 home_ss.dll
68d80000 00050000 hnetwiz.dll
68de0000 00010000 hnetmon.dll
68df0000 00040000 hnetcfg.dll
68e40000 00010000 hmmapi.dll
68e50000 00010000 hidserv.dll
68e60000 00010000 hid.dll
68e70000 00020000 hhctrlui.dll
68e90000 00010000 hexedit.dll
68ea0000 00010000 hcappres.dll
68eb0000 000a0000 h323msp.dll
68f50000 00010000 gzip.dll
68f60000 00030000 guitrn_a.dll
68f90000 00030000 guitrn.dll
68fc0000 00010000 grovmsg.dll
68fd0000 00030000 gptext.dll
69000000 00010000 gpkrsrc.dll
69010000 00080000 gpedit.dll
69090000 00020000 glu32.dll
690c0000 00050000 glmf32.dll
69110000 000a0000 getuname.dll
691b0000 00020000 gcdef.dll
691d0000 00070000 fxsxp32.dll
69240000 00030000 fxswzrd.dll
69280000 00030000 fxsui.dll
692b0000 00070000 fxstiff.dll
69320000 00010000 fxst30p.dll
69330000 00040000 fxst30.dll
69370000 00090000 fxsst.dll
69400000 00020000 fxsrtmtd.dll
69420000 00010000 fxsroute.dll
69430000 00010000 fxsres.dll
69440000 00010000 fxsperf.dll
69450000 00030000 fxsocm.dll
69480000 00010000 fxsmon.dll
69490000 00010000 fxsext32.dll
694a0000 00020000 fxsevent.dll
694c0000 00010000 fxsdrv.dll
694d0000 00050000 fxscomex.dll
69520000 00020000 fxscom.dll
69540000 00030000 fxsclntr.dll
69570000 00020000 fxscfgwz.dll
69590000 00070000 fxsapi.dll
69610000 00070000 fxsadmin.dll
69680000 00010000 fx5eres.dll
69690000 00020000 fwdprov.dll
696b0000 00020000 fuusd.dll
696d0000 00030000 fupclres.dll
69700000 00010000 fu9res.dll
69710000 00010000 fu24res.dll
69720000 00030000 ftsrch.dll
69760000 00020000 ftpsvc2.dll
69790000 00020000 ftpsv251.dll
697c0000 00010000 ftpsapi2.dll
697d0000 00010000 ftpmib.dll
697e0000 00010000 ftpctrs2.dll
697f0000 00010000 ftlx041e.dll
69800000 00020000 fsusd.dll
69820000 00010000 fsconins.dll
69830000 00010000 fscfg.dll
69840000 00030000 framedyn.dll
69870000 00010000 fpnwclnt.dll
69880000 00010000 fp40ext.dll
69890000 00020000 fontsub.dll
698b0000 00060000 fontext.dll
69920000 00020000 fnfilter.dll
69940000 00010000 fmifs.dll
69950000 00020000 fldrclnr.dll
69970000 00010000 feclient.dll
69980000 00020000 fdeploy.dll
699a0000 00030000 fde.dll
699d0000 00020000 faultrep.dll
699f0000 00010000 f3ahvoas.dll
69a00000 00030000 exts.dll
69a30000 00010000 exstrace.dll
69a40000 00010000 exp24res.dll
69a50000 00010000 evtgprov.dll
69a60000 00010000 evntrprv.dll
69a70000 00020000 evntagnt.dll
69a90000 00010000 eventcls.dll
69aa0000 00010000 pidgen.dll
69ab0000 00010000 esunid.dll
69ad0000 00010000 esunib.dll
69af0000 00010000 esuni.dll
69b10000 00020000 esuimgd.dll
69b30000 00010000 esuimg.dll
69b40000 00010000 esucmd.dll
69b50000 00010000 esucm.dll
69b60000 00010000 esentprf.dll
69b70000 00120000 esent97.dll
69c90000 00100000 esent.dll
69d90000 00010000 escp2res.dll
69da0000 00010000 es1371mp.dll
69db0000 00020000 eqnclass.dll
69dd0000 00010000 epnutx22.dll
69de0000 00120000 epnhtx2h.dll
69f00000 00090000 epnhtx16.dll
69f90000 000a0000 epnhtx15.dll
6a030000 00090000 epnhtx14.dll
6a0d0000 00090000 epnhtx13.dll
6a160000 00080000 epnhtx12.dll
6a1e0000 00090000 epnhtx11.dll
6a270000 00060000 epnhtx0a.dll
6a2d0000 00060000 epnhtx09.dll
6a330000 00070000 epnhtx07.dll
6a3a0000 00070000 epnhtx05.dll
6a410000 00060000 epnhtx04.dll
6a470000 00060000 epnhtx02.dll
6a4d0000 00060000 epnhtx01.dll
6a530000 00160000 epnhte5d.dll
6a690000 00140000 epnhte5a.dll
6a7d0000 00140000 epnhte4s.dll
6a910000 00110000 epnhte4p.dll
6aa20000 00190000 epnhte4n.dll
6abb0000 00170000 epnhte4l.dll
6ad20000 00220000 epnhte4k.dll
6af40000 00200000 epnhte4j.dll
6b140000 00140000 epnhte4i.dll
6b280000 00130000 epnhte4h.dll
6b3b0000 00130000 epnhte4g.dll
6b4e0000 00090000 epnhte4d.dll
6b570000 00110000 epnhte4c.dll
6b680000 00110000 epnhte4b.dll
6b790000 000b0000 epnhte4a.dll
6b840000 000f0000 epnhte3v.dll
6b930000 001b0000 epnhte3t.dll
6bae0000 00160000 epnhte3q.dll
6bc40000 00060000 epnhte3p.dll
6bca0000 00070000 epnhte3o.dll
6bd10000 000f0000 epnhte3n.dll
6be00000 000a0000 epnhte2m.dll
6bea0000 000e0000 epnhte2k.dll
6bf80000 00140000 epnhte2j.dll
6c0c0000 00020000 epngui40.dll
6c0e0000 00020000 epngui30.dll
6c100000 00020000 epngui10.dll
6c120000 00010000 epndrv01.dll
6c130000 00020000 eplvcd00.dll
6c150000 00020000 eplrcz00.dll
6c170000 00010000 epcl5ui.dll
6c180000 00020000 epcl5res.dll
6c1b0000 00010000 ep9res.dll
6c1c0000 00010000 ep9bres.dll
6c1d0000 00020000 ep2bres.dll
6c1f0000 00010000 ep24res.dll
6c200000 00010000 efsadu.dll
6c210000 00110000 edb500.dll
6c330000 00010000 ecp2eres.dll
6c350000 00040000 dxtrans.dll
6c390000 00060000 dxtmsft.dll
6c3f0000 000e0000 dxmrtp.dll
6c4d0000 00080000 dxmasf.dll
6c550000 00130000 dx8vb.dll
6c680000 000a0000 dx7vb.dll
6c720000 00010000 dvusd.dll
6c730000 00050000 duser.dll
6c780000 00010000 dswave.dll
6c790000 00020000 dsuiwiz.dll
6c7b0000 00020000 dsuiext.dll
6c7d0000 00010000 dssec.dll
6c7e0000 00040000 dsquery.dll
6c820000 00020000 dsprov.dll
6c850000 00030000 dsprop.dll
6c880000 00140000 dsound3d.dll
6c9d0000 00030000 dskquoui.dll
6ca00000 00020000 dskquota.dll
6ca20000 00020000 dsdmoprp.dll
6ca40000 00030000 dsdmo.dll
6ca70000 00020000 dsauth.dll
6ca90000 00090000 dsadmin.dll
6cb30000 00020000 drmstor.dll
6cb50000 00010000 dpwsockx.dll
6cb70000 00010000 dpwsock.dll
6cb80000 00020000 dpvvox.dll
6cba0000 00040000 dpvoice.dll
6cbe0000 00010000 dpvacm.dll
6cbf0000 00010000 dpserial.dll
6cc10000 00020000 dpnwsock.dll
6cc30000 00020000 dpnmodem.dll
6cc50000 00010000 dpnlobby.dll
6cc60000 00020000 dpnhupnp.dll
6cc80000 00010000 dpnhpast.dll
6cc90000 00030000 dpnet.dll
6ccc0000 00010000 dpnaddr.dll
6ccd0000 00010000 dpmodemx.dll
6cce0000 00040000 dplayx.dll
6cd20000 00020000 dplay.dll
6cd40000 00040000 dpcres.dll
6cd80000 00020000 dpcdll.dll
6cdb0000 00020000 domadmin.dll
6cdd0000 00010000 docprop2.dll
6cde0000 00010000 docprop.dll
6ce00000 00030000 dnsprov.dll
6ce30000 00010000 dnsperf.dll
6ce40000 000d0000 dnsmgr.dll
6cf10000 00020000 dmusic.dll
6cf30000 00020000 dmsynth.dll
6cf50000 00020000 dmstyle.dll
6cf70000 00020000 dmscript.dll
6cf90000 00010000 dmocx.dll
6cfa0000 00010000 dmloader.dll
6cfb0000 00010000 dmintf.dll
6cfc0000 00030000 dmime.dll
6d000000 00050000 dmdlgs.dll
6d050000 000d0000 dmconfig.dll
6d130000 00020000 dmcompos.dll
6d150000 00010000 dmband.dll
6d160000 00020000 divasu.dll
6d180000 00020000 divaprop.dll
6d1a0000 00010000 divaci.dll
6d1b0000 00020000 disrvsu.dll
6d1d0000 00010000 disrvpp.dll
6d1e0000 00010000 disrvci.dll
6d1f0000 00010000 dispex.dll
6d200000 00180000 diskcopy.dll
6d380000 00020000 directdb.dll
6d3a0000 00040000 dinput8.dll
6d3e0000 00010000 dimap.dll
6d3f0000 00020000 digirlpt.dll
6d410000 00010000 digiisdn.dll
6d420000 00020000 digiinf.dll
6d440000 00030000 digihlc.dll
6d470000 00040000 digifwrk.dll
6d4b0000 00020000 digidbp.dll
6d4e0000 00010000 digiasyn.dll
6d500000 00010000 diconres.dll
6d510000 00010000 diapi2nt.dll
6d520000 00010000 diapi232.dll
6d530000 00070000 diactfrm.dll
6d5a0000 00050000 dhcpssvc.dll
6d5f0000 000f0000 dhcpsnap.dll
6d6e0000 00020000 dhcpsapi.dll
6d700000 00070000 dhcpmon.dll
6d770000 00010000 dhcpmib.dll
6d780000 00020000 dgsetup.dll
6d7a0000 00030000 dgrpsetu.dll
6d7d0000 00030000 dgnet.dll
6d800000 00070000 dgconfig.dll
6d870000 00010000 dgclass.dll
6d880000 00010000 dfsshlex.dll
6d890000 00010000 dfssetup.dll
6d8a0000 00060000 dfsgui.dll
6d900000 00020000 dfscore.dll
6d920000 00030000 dfrgui.dll
6d950000 00010000 dfrgsnap.dll
6d960000 00010000 dfrgres.dll
6d980000 00010000 deskperf.dll
6d990000 00010000 deskmon.dll
6d9a0000 00010000 deskadp.dll
6d9b0000 00010000 debugex.dll
6d9c0000 00010000 ddrawex.dll
6d9d0000 00010000 dcpromo.dll
6d9e0000 00010000 dclsres.dll
6d9f0000 00010000 dc9res.dll
6da00000 00020000 dc260usd.dll
6da20000 00010000 dc24res.dll
6da30000 00020000 dc240usd.dll
6da50000 00020000 dc210usd.dll
6da70000 00010000 dc210_32.dll
6da80000 00020000 dbnetlib.dll
6daa0000 00080000 dbghelp.dll
6db20000 00100000 dbgeng.dll
6dc20000 00030000 datime.dll
6dc50000 00010000 dataclen.dll
6dc70000 00100000 danim.dll
6dd70000 00020000 d3dxof.dll
6dd90000 00060000 d3drm.dll
6ddf0000 000a0000 d3dramp.dll
6de90000 00010000 d3dpmesh.dll
6dea0000 00080000 d3dim.dll
6df20000 00010000 d3d8thk.dll
6df30000 00130000 d3d8.dll
6e060000 00010000 cyzports.dll
6e070000 00010000 cyzcoins.dll
6e080000 00010000 cyyports.dll
6e090000 00010000 cyycoins.dll
6e0a0000 00010000 ctmrclas.dll
6e0b0000 00040000 ctmasetp.dll
6e0f0000 00020000 ctl3d32.dll
6e110000 00010000 ct9res.dll
6e120000 00020000 ct24res.dll
6e140000 00020000 csseqchk.dll
6e160000 00010000 csapi3t1.dll
6e180000 00030000 csamsp.dll
6e1b0000 00010000 cryptext.dll
6e1c0000 00020000 cryptdlg.dll
6e1e0000 000f0000 cqsdclr2.dll
6e2d0000 001c0000 cqsdclr1.dll
6e490000 00030000 cq90sui.dll
6e4c0000 00010000 cq90sres.dll
6e4d0000 00010000 cq90srdr.dll
6e4e0000 00060000 cq90icur.dll
6e540000 00020000 cq90fcic.dll
6e570000 00030000 cq75sui.dll
6e5a0000 00010000 cq75sres.dll
6e5b0000 00010000 cq75srdr.dll
6e5c0000 00060000 cq75icur.dll
6e620000 00030000 cq75fcic.dll
6e650000 00030000 cq70sui.dll
6e680000 00010000 cq70sres.dll
6e690000 00010000 cq70srdr.dll
6e6a0000 00060000 cq70icur.dll
6e700000 00020000 cq70fcic.dll
6e730000 00030000 cq60sui.dll
6e760000 00010000 cq60sres.dll
6e770000 00010000 cq60srdr.dll
6e780000 00060000 cq60icur.dll
6e7e0000 00030000 cq60fcic.dll
6e810000 00030000 cq30sui.dll
6e840000 00010000 cq30sres.dll
6e850000 00010000 cq30srdr.dll
6e860000 00060000 cq30icur.dll
6e8c0000 00030000 cq30fcic.dll
6e8f0000 00030000 cq12sui.dll
6e920000 00010000 cq12sres.dll
6e930000 00010000 cq12srdr.dll
6e940000 00060000 cq12icur.dll
6e9a0000 00030000 cq12fcic.dll
6e9d0000 00050000 cpscan.dll
6ea20000 00010000 counters.dll
6ea30000 00010000 corpol.dll
6ea40000 00010000 convmsg.dll
6ea50000 00010000 controt.dll
6ea60000 00020000 console.dll
6ea80000 00060000 confmsp.dll
6eae0000 00010000 confmrsl.dll
6eaf0000 00080000 comuid.dll
6eb70000 00030000 comsnap.dll
6eba0000 00050000 comsetup.dll
6ebf0000 00020000 comrepl.dll
6ec10000 00040000 compstui.dll
6ec50000 00010000 compfilt.dll
6ec60000 00040000 compatui.dll
6ecb0000 00010000 comcat.dll
6ecc0000 00040000 comadmin.dll
6ed00000 00010000 comaddin.dll
6ed10000 00010000 coadmin.dll
6ed20000 00010000 cnvfat.dll
6ed30000 00010000 cnusd.dll
6ed40000 00020000 cnlbpres.dll
6ed60000 00010000 cnetcfg.dll
6ed70000 00010000 cnbs4500.dll
6ed80000 00010000 cnbs450.dll
6ed90000 00010000 cnbs400.dll
6eda0000 00010000 cnbpgr08.dll
6edb0000 00030000 cnbpgr05.dll
6ede0000 00040000 cnbpgr03.dll
6ee20000 00010000 cnbpgr02.dll
6ee30000 00010000 cnbpgr01.dll
6ee40000 00010000 cnbostd.dll
6ee50000 00010000 cnbo64.dll
6ee60000 00010000 cnbo59.dll
6ee70000 00050000 cnbjui2.dll
6eec0000 00040000 cnbjui.dll
6ef00000 00020000 cnbjmon2.dll
6ef20000 00020000 cnbjdrv2.dll
6ef40000 00020000 cnbjdrv.dll
6ef60000 00020000 cnbjdrs.dll
6ef80000 00070000 cnbjdrc.dll
6eff0000 00010000 cnbjcres.dll
6f000000 00010000 cnb85.dll
6f010000 00010000 cnb820.dll
6f020000 00010000 cnb8000.dll
6f030000 00010000 cnb800.dll
6f040000 00010000 cnb80.dll
6f050000 00010000 cnb7100.dll
6f060000 00010000 cnb7000.dll
6f070000 00010000 cnb70.dll
6f080000 00010000 cnb6500.dll
6f090000 00010000 cnb6200.dll
6f0a0000 00010000 cnb620.dll
6f0b0000 00010000 cnb6100.dll
6f0c0000 00010000 cnb610.dll
6f0d0000 00010000 cnb600e.dll
6f0e0000 00010000 cnb6000.dll
6f0f0000 00010000 cnb600.dll
6f100000 00010000 cnb5500.dll
6f110000 00010000 cnb55.dll
6f120000 00010000 cnb50.dll
6f130000 00010000 cnb4650.dll
6f140000 00010000 cnb4550.dll
6f150000 00010000 cnb4400.dll
6f160000 00010000 cnb4300s.dll
6f170000 00010000 cnb4300.dll
6f180000 00010000 cnb4200s.dll
6f190000 00010000 cnb4200.dll
6f1a0000 00010000 cnb4100.dll
6f1b0000 00010000 cnb4000.dll
6f1c0000 00010000 cnb3000.dll
6f1d0000 00010000 cnb265sp.dll
6f1e0000 00010000 cnb255sp.dll
6f1f0000 00010000 cnb250.dll
6f200000 00010000 cnb240.dll
6f210000 00010000 cnb210sp.dll
6f220000 00010000 cnb2100s.dll
6f230000 00010000 cnb2100.dll
6f240000 00010000 cnb210.dll
6f250000 00010000 cnb2000s.dll
6f260000 00010000 cnb2000.dll
6f270000 00010000 cnb1000s.dll
6f280000 00010000 cnb1000.dll
6f290000 00010000 cn330res.dll
6f2a0000 00010000 cn32602.dll
6f2b0000 00010000 cn32601.dll
6f2c0000 00010000 cn32600.dll
6f2e0000 00010000 cn2002.dll
6f2f0000 00020000 cn2001.dll
6f310000 00010000 cn2000.dll
6f330000 00010000 cn1760e2.dll
6f340000 00010000 cn1760e1.dll
6f350000 00020000 cn1760e0.dll
6f370000 00010000 cn1602.dll
6f380000 00010000 cn1601.dll
6f390000 00010000 cn1600.dll
6f3b0000 00010000 cn10002.dll
6f3c0000 00010000 cn10001.dll
6f3d0000 00010000 cn10000.dll
6f3f0000 00020000 cmutoa.dll
6f410000 00010000 cmutil.dll
6f420000 00010000 cmroute.dll
6f430000 00010000 cmproxy.dll
6f440000 00040000 cmprops.dll
6f480000 00010000 cmpbk32.dll
6f490000 00110000 cmnresm.dll
6f5a0000 00040000 cmnclim.dll
6f5e0000 00060000 cmdial32.dll
6f640000 00010000 cmcfg32.dll
6f650000 00020000 cluswmi.dll
6f670000 00010000 clussprt.dll
6f680000 00060000 clusres.dll
6f6e0000 00010000 clusocm.dll
6f6f0000 00010000 clusiis4.dll
6f700000 00010000 cluadmmc.dll
6f720000 00030000 cluadmex.dll
6f750000 00010000 clnetrex.dll
6f770000 00010000 clnetres.dll
6f780000 00090000 clcfgsrv.dll
6f820000 00020000 clbcatex.dll
6f840000 00010000 clb.dll
6f850000 00070000 class_ss.dll
6f8c0000 00050000 cladmwiz.dll
6f910000 00010000 citohres.dll
6f920000 00020000 ciodm.dll
6f940000 00140000 cimwin32.dll
6fa80000 00020000 cic.dll
6faa0000 00030000 ciadmin.dll
6fad0000 000d0000 chkrres.dll
6fba0000 00010000 chkr.dll
6fbb0000 00010000 cfgbkend.dll
6fbc0000 00030000 cewmdm.dll
6fc00000 00010000 certxds.dll
6fc10000 00040000 certtmpl.dll
6fc50000 00020000 certpdef.dll
6fc70000 00040000 certocm.dll
6fcc0000 00020000 certobj.dll
6fce0000 00070000 certmmc.dll
6fd50000 00080000 certmgr.dll
6fdd0000 00010000 certenc.dll
6fde0000 00020000 certdb.dll
6fe00000 00020000 certadm.dll
6fe20000 001f0000 cdosys.dll
70020000 00010000 cdmodem.dll
70030000 00010000 cdm.dll
70040000 00030000 cdfview.dll
70070000 00010000 ccfgnt.dll
70080000 00010000 ccfg95.dll
70090000 00020000 ccfapi32.dll
700b0000 000a0000 catsrvut.dll
70150000 00020000 catsrvps.dll
70170000 00040000 catsrv.dll
701b0000 00060000 cards.dll
70210000 00030000 capesnpn.dll
70240000 00010000 camocx.dll
70250000 00020000 camext30.dll
70280000 00040000 camext20.dll
702c0000 00020000 camexo20.dll
702e0000 00020000 cabview.dll
70300000 00010000 c_iscii.dll
70310000 00010000 c_is2022.dll
70320000 00040000 c_g18030.dll
70360000 00010000 bull9res.dll
70380000 00020000 bul24res.dll
703a0000 00010000 bul18res.dll
703b0000 00010000 btpagnt.dll
703c0000 00010000 brserif.dll
703d0000 00010000 brscnrsm.dll
703e0000 00010000 brpinfo.dll
703f0000 00020000 browsewm.dll
70410000 00010000 browscap.dll
70420000 00010000 brothui.dll
70430000 00010000 brother.dll
70440000 00020000 brmfusb.dll
70460000 00010000 brmfpmon.dll
70470000 00030000 brmflpt.dll
704a0000 00020000 brmfcwia.dll
704c0000 00010000 brmfbidi.dll
704d0000 000a0000 brhlres.dll
70570000 00010000 brhjres.dll
70580000 00010000 brevif.dll
70590000 00020000 brcoinst.dll
705b0000 00010000 brclrui.dll
705c0000 00010000 brclr0ui.dll
705d0000 000f0000 brclr00.dll
706c0000 00080000 brclr0.dll
70740000 00080000 brclr.dll
707c0000 00010000 brcl00ui.dll
707d0000 00010000 brbidiif.dll
707e0000 00010000 br9res.dll
707f0000 00010000 br24res.dll
70810000 00030000 bnts.dll
70840000 00060000 blue_ss.dll
708a0000 00020000 binlsvc.dll
708c0000 00010000 bidispl.dll
708d0000 00010000 bhsupp.dll
708e0000 00010000 bhp025.dll
708f0000 00010000 bhp024.dll
70900000 00010000 bhp023.dll
70910000 00010000 bhp022.dll
70920000 00020000 bhp021.dll
70950000 00020000 bhp020.dll
70970000 00030000 bhp019.dll
709a0000 00010000 bhp018.dll
709b0000 00010000 bhp017.dll
709c0000 00010000 bhp016.dll
709d0000 00040000 bhp015.dll
70a10000 00010000 bhp014.dll
70a20000 00030000 bhp013.dll
70a50000 00010000 bhp012.dll
70a60000 00010000 bhp011.dll
70a70000 00010000 bhp010.dll
70a80000 00030000 bhp009.dll
70ab0000 00010000 bhp008.dll
70ac0000 00020000 bhp007.dll
70ae0000 00010000 bhp006.dll
70af0000 00010000 bhp005.dll
70b00000 00010000 bhp004.dll
70b10000 00010000 bhp003.dll
70b20000 00010000 bhp002.dll
70b30000 00020000 bhp001.dll
70b50000 001c0000 bckgres.dll
70d20000 00020000 bckg.dll
70d40000 00010000 batt.dll
70d50000 00020000 avwav.dll
70d70000 00040000 avtapi.dll
70db0000 00010000 avmeter.dll
70dc0000 00030000 avmenum.dll
70df0000 00020000 avmcoxp.dll
70e10000 00010000 avmc2032.dll
70e20000 00020000 autodisc.dll
70e40000 00010000 authfilt.dll
70e50000 00010000 audiosrv.dll
70e60000 00010000 atrace.dll
70e70000 00010000 atmpvcno.dll
70e80000 00010000 atkctrs.dll
70e90000 00020000 asycfilt.dll
70eb0000 00010000 asptxn.dll
70ec0000 00010000 aspperf.dll
70ed0000 00060000 asp51.dll
70f30000 00060000 asp.dll
70f90000 00010000 asfsipc.dll
70fa0000 00010000 asferror.dll
70fb0000 00050000 appmgr.dll
71000000 00020000 appconf.dll
71020000 00020000 apcups.dll
71040000 00020000 amstream.dll
71060000 00010000 alrsvc.dll
71070000 00010000 alpsres.dll
71090000 00030000 air300pp.dll
710c0000 00010000 agtintl.dll
710d0000 00010000 agt0c0a.dll
710e0000 00010000 agt0816.dll
710f0000 00010000 agt0804.dll
71100000 00010000 agt041f.dll
71110000 00010000 agt041d.dll
71120000 00010000 agt0419.dll
71130000 00010000 agt0416.dll
71140000 00010000 agt0415.dll
71150000 00010000 agt0414.dll
71160000 00010000 agt0413.dll
71170000 00010000 agt0412.dll
71180000 00010000 agt0411.dll
71190000 00010000 agt0410.dll
711a0000 00010000 agt040e.dll
711b0000 00010000 agt040d.dll
711c0000 00010000 agt040c.dll
711d0000 00010000 agt040b.dll
711e0000 00010000 agt0409.dll
711f0000 00010000 agt0408.dll
71200000 00010000 agt0407.dll
71210000 00010000 agt0406.dll
71220000 00010000 agt0405.dll
71230000 00010000 agt0404.dll
71240000 00010000 agt0401.dll
71250000 00010000 agentsr.dll
71260000 00010000 agentpsh.dll
71270000 00010000 agentmpx.dll
71280000 00010000 agentdpv.dll
712a0000 00010000 agentdp2.dll
712b0000 00040000 agentctl.dll
712f0000 00010000 agentanm.dll
71300000 00020000 adsnw.dll
71320000 00030000 adsnds.dll
71350000 00020000 adsmsext.dll
71370000 00030000 adsldp.dll
713a0000 00050000 adsiis51.dll
713f0000 00050000 adsiis.dll
71440000 00010000 adrot.dll
71460000 000b0000 adprop.dll
71510000 00010000 admxprox.dll
71520000 00010000 admwprox.dll
71530000 00020000 admparse.dll
71550000 00010000 admexs.dll
71560000 00020000 acxtrnal.dll
71590000 00030000 input.dll
715c0000 00070000 acspecfc.dll
71630000 00020000 aclui.dll
71650000 00010000 OPEN
71670000 00080000 aclayers.dll
716f0000 00030000 aclua.dll
71720000 00050000 acverfyr.dll
71770000 000b0000 appwiz.cpl
71820000 00020000 OPEN
71840000 00020000 acerscad.dll
71860000 00020000 acctres.dll
71880000 00010000 aaaamon.dll
71890000 00080000 a3dapi.dll
71910000 00030000 a3d.dll
71940000 00010000 OPEN
71950000 00030000 31x5us04.dll
71980000 00030000 31x5uc04.dll
719b0000 00030000 31x5rs04.dll
719e0000 00030000 31x5rc04.dll
71a10000 00010000 31x5ls04.dll
71a20000 00010000 31x5lc04.dll
71a30000 00010000 msafd.dll
71a40000 00040000 mswsock.dll
71a80000 00010000 wshtcpip.dll
71a90000 00010000 ws2help.dll
71aa0000 00020000 ws2_32.dll
71ac0000 00010000 wsock32.dll
71ad0000 00020000 ntlanui.dll
71af0000 00010000 mprui.dll
71b10000 00020000 mpr.dll
71b30000 00030000 netmsg.dll
71b60000 00030000 acledit.dll
71b90000 00050000 netui2.dll
71be0000 00020000 samlib.dll
71c00000 00010000 ntlanman.dll
71c10000 00050000 netapi32.dll
71c70000 00010000 netrap.dll
71c80000 00040000 netui1.dll
71cc0000 00020000 netui0.dll
71ce0000 00050000 kerberos.dll
71d30000 00020000 actxprxy.dll
71d50000 00030000 msconv97.dll
71d80000 00020000 url.dll
71da0000 00040000 syncui.dll
71de0000 00010000 olesvr32.dll
71df0000 00010000 olecnv32.dll
71e00000 00020000 olecli32.dll
71e20000 00020000 olethk32.dll
71e40000 00020000 msapsspc.dll
71e60000 00020000 6to4svc.dll
71e80000 00010000 OPEN
71e90000 00010000 ntdsbcli.dll
71ea0000 00010000 ntdsbsrv.dll
71eb0000 00020000 ntdsetup.dll
71ed0000 00010000 hticons.dll
71ee0000 00040000 netevent.dll
71f20000 00010000 wshisn.dll
71f30000 00010000 w32topl.dll
71f40000 00010000 wshnetbs.dll
71f50000 00010000 snmpapi.dll
71f60000 00010000 ipxwan.dll
71f70000 00010000 security.dll
71f80000 00010000 ureg.dll
71f90000 00050000 ulib.dll
71fe0000 00010000 ntdsatq.dll
71ff0000 00010000 uniplat.dll
72000000 00010000 wsnmp32.dll
72010000 00010000 mgmtapi.dll
72020000 00010000 tcpmib.dll
72030000 00020000 adptif.dll
72050000 00010000 rastapi.dll
72070000 00020000 xactsrv.dll
72090000 00020000 rasauto.dll
720b0000 00020000 ntdskcc.dll
720d0000 00010000 mssign32.dll
720e0000 00150000 ntdsa.dll
72230000 00040000 rasppp.dll
72270000 00030000 dinput.dll
722a0000 00010000 sensapi.dll
722b0000 00010000 winfax.dll
722c0000 00010000 sens.dll
722d0000 00070000 ntmssvc.dll
72340000 00030000 ntmsdba.dll
72370000 00020000 polstore.dll
72390000 00010000 mmcshext.dll
723a0000 00020000 hhsetup.dll
723c0000 00020000 winscard.dll
723e0000 00010000 usbmon.dll
723f0000 00010000 tcpmon.dll
72400000 00020000 mydocs.dll
72420000 00020000 browselc.dll
72440000 00010000 rnr20.dll
72450000 00030000 rasmans.dll
72480000 00010000 ntlsapi.dll
72490000 00010000 mspmspsv.dll
724b0000 00060000 smlogcfg.dll
72510000 00010000 rassapi.dll
72520000 00050000 pdh.dll
72580000 00080000 ntmsmgr.dll
72600000 00010000 ntmsapi.dll
72610000 00020000 mycomput.dll
72630000 00080000 msxml.dll
726c0000 00120000 mmcndmgr.dll
727e0000 00020000 mmcbase.dll
72800000 00100000 mfc42u.dll
72900000 00040000 localsec.dll
72940000 00060000 filemgmt.dll
729a0000 00030000 els.dll
729d0000 00010000 dmutil.dll
729f0000 00030000 dmdskres.dll
72a20000 00030000 dmdskmgr.dll
72a60000 00050000 devmgr.dll
72ab0000 00040000 adsnt.dll
72af0000 00020000 plugin.ocx
72b10000 000a0000 mstscax.dll
72bb0000 00010000 xrxnps.dll
72bc0000 000e0000 msdxm.ocx
72ca0000 00020000 l3codecx.ax
72cc0000 00010000 msadp32.acm
72cd0000 00010000 zeeverm.dll
72ce0000 00010000 msacm32.drv
72cf0000 00010000 wdmaud.drv
72d00000 000d0000 xxui1.dll
72dd0000 00120000 msxml3.dll
72ef0000 00030000 wmiprov.dll
72f20000 00010000 zoneoc.dll
72f30000 00020000 loadperf.dll
72f50000 00020000 wmimsg.dll
72f70000 00060000 usp10.dll
72fd0000 00030000 winspool.drv
73000000 00010000 wzcsapi.dll
73010000 00010000 rrcm.dll
73020000 00010000 nmasnt.dll
73030000 00010000 h323cc.dll
73040000 00010000 dcap32.dll
73050000 00020000 rsvpsp.dll
73070000 00020000 nmcom.dll
73090000 00020000 nmchat.dll
730b0000 00040000 nmas.dll
730f0000 00040000 nac.dll
73130000 00040000 mst120.dll
73170000 00060000 callcont.dll
731d0000 000c0000 winntbba.dll
732a0000 00010000 softpub.dll
732b0000 00010000 riched32.dll
732c0000 00010000 mscat32.dll
732d0000 00080000 vbscript.dll
73350000 00060000 zipfldr.dll
733b0000 00040000 tapisrv.dll
733f0000 00160000 msvbvm60.dll
73550000 00010000 zonelibm.dll
73560000 00010000 traffic.dll
73570000 00030000 scrrun.dll
735a0000 00040000 mstask.dll
735f0000 00010000 digest.dll
73610000 00010000 mnmdd.dll
73620000 00020000 mciavi32.dll
73640000 00010000 tsbyuv.dll
73650000 00010000 msyuv.dll
73660000 00010000 msvidc32.dll
73670000 00010000 msrle32.dll
73680000 00010000 msdmo.dll
73690000 00010000 iyuv_32.dll
736a0000 00030000 qcap.dll
736e0000 00050000 ir50_qcx.dll
73730000 00050000 ddraw.dll
73780000 00060000 ir41_qcx.dll
737e0000 00060000 ir32_32.dll
73840000 000d0000 ir50_32.dll
73910000 000d0000 d3dim700.dll
739e0000 00020000 xrxwiadr.dll
73a10000 00060000 wiaservc.dll
73a70000 00010000 znetm.dll
73a80000 00020000 zoneclim.dll
73ab0000 00050000 msvcrt20.dll
73b00000 00020000 mscms.dll
73b20000 00020000 avifil32.dll
73b40000 00010000 tsd32.dll
73b50000 00020000 avicap32.dll
73b70000 00020000 sti.dll
73b90000 00010000 dciman32.dll
73ba0000 00020000 msvfw32.dll
73bd0000 00020000 iccvid.dll
73bf0000 00010000 atmlib.dll
73c00000 000b0000 spxports.dll
73cb0000 00040000 t2embed.dll
73cf0000 00010000 seclogon.dll
73d00000 00020000 wbemcons.dll
73d20000 00010000 cryptnet.dll
73d40000 00020000 shgina.dll
73d60000 00030000 crtdll.dll
73d90000 00010000 lz32.dll
73da0000 00100000 mfc42.dll
73ea0000 00010000 mmdrv.dll
73eb0000 00010000 ksuser.dll
73ec0000 00010000 devenum.dll
73ee0000 00060000 dsound.dll
73f40000 00150000 quartz.dll
74090000 00150000 msvbvm50.dll
741e0000 00020000 sfman32.dll
74200000 00050000 devcon32.dll
74250000 00010000 pjlmon.dll
74260000 00010000 icmp.dll
74270000 00010000 cnbjmon.dll
74280000 00020000 win32spl.dll
742b0000 00020000 spoolss.dll
742d0000 00020000 inetpp.dll
742f0000 00050000 localspl.dll
74340000 00010000 winipsec.dll
74350000 00010000 wdigest.dll
74370000 00010000 pstorsvc.dll
74380000 00010000 msprivs.dll
74390000 00020000 psbase.dll
743b0000 00030000 ipsecsvc.dll
743e0000 00030000 scecli.dll
74410000 00070000 samsrv.dll
74480000 00070000 netlogon.dll
744f0000 000b0000 lsasrv.dll
745a0000 000c0000 oakley.dll
74660000 00030000 xuim760.dll
74690000 00030000 msls31.dll
746c0000 00030000 msimtf.dll
746f0000 00050000 msctf.dll
74740000 00090000 mlang.dll
747e0000 002c0000 mshtml.dll
74aa0000 00010000 powrprof.dll
74ab0000 00010000 cfgmgr32.dll
74ac0000 00010000 batmeter.dll
74ad0000 00020000 stobject.dll
74b00000 00050000 webcheck.dll
74b50000 00090000 printui.dll
74be0000 00010000 ssdpsrv.dll
74bf0000 00010000 regsvc.dll
74c10000 00010000 lmhsvc.dll
74c20000 00020000 msdart.dll
74c50000 00030000 oleacc.dll
74c80000 00070000 mshtmled.dll
74d00000 00020000 oledlg.dll
74d30000 00020000 msoert2.dll
74d60000 000a0000 inetcomm.dll
74e00000 00070000 riched20.dll
74e70000 00010000 wshext.dll
74e90000 00010000 wuauserv.dll
74ea0000 00010000 wbemsvc.dll
74ec0000 00010000 wbemprox.dll
74ed0000 00010000 ssdpapi.dll
74ee0000 00020000 rastls.dll
74f00000 00010000 xxpsru1.dll
74f10000 00010000 pchsvc.dll
74f20000 00010000 msidle.dll
74f30000 00010000 msgsvc.dll
74f40000 00010000 icaapi.dll
74f50000 00010000 ersvc.dll
74f60000 00010000 dmserver.dll
74f70000 00010000 cryptsvc.dll
74f90000 00020000 clusapi.dll
74fb0000 00010000 browser.dll
74fd0000 00020000 raschap
74ff0000 00020000 wmiutils.dll
75010000 00030000 upnp.dll
75040000 00020000 trkwks.dll
75060000 00020000 srvsvc.dll
75080000 00020000 resutils.dll
750a0000 00020000 mtxoci.dll
750c0000 00020000 mtxclu.dll
750e0000 00020000 mstlsapi.dll
75100000 00020000 colbact.dll
75120000 00020000 cabinet.dll
75140000 00020000 wkssvc.dll
75170000 00030000 srsvc.dll
751a0000 00030000 schedsvc.dll
751d0000 00030000 repdrvfs.dll
75200000 00030000 appmgmts.dll
75230000 00030000 advpack.dll
75260000 00040000 wbemcomn.dll
752a0000 00040000 termsrv.dll
752e0000 00040000 esscli.dll
75320000 00040000 certcli.dll
75360000 00050000 wbemess.dll
753b0000 00070000 vssapi.dll
75420000 00080000 wbemcore.dll
754a0000 00080000 cryptui.dll
75520000 000a0000 rasdlg.dll
755d0000 000a0000 netcfgx.dll
75670000 000a0000 fastprox.dll
75710000 00120000 comsvcs.dll
75830000 00050000 rpcss.dll
75880000 00010000 eventlog.dll
758a0000 00020000 umpnpmgr.dll
758c0000 00050000 scesrv.dll
75910000 00010000 profmap.dll
75920000 00010000 nddeapi.dll
75930000 00020000 wlnotify.dll
75950000 00100000 msgina.dll
75a50000 000b0000 userenv.dll
75b00000 00020000 xcci2032.dll
75b20000 00010000 csrsrv.dll
75b30000 00010000 basesrv.dll
75b40000 00050000 winsrv.dll
75b90000 000a0000 unires.dll
75c30000 000a0000 jscript.dll
75cd0000 001a0000 netshell.dll
75e70000 000b0000 sxs.dll
75f20000 00020000 apphelp.dll
75f40000 00010000 drprov.dll
75f50000 00010000 davclnt.dll
75f60000 00100000 browseui.dll
76060000 00070000 msvcp60.dll
760d0000 00080000 urlmon.dll
76150000 00090000 shdoclc.dll
761e0000 000a0000 wininet.dll
76280000 00010000 msasn1.dll
762a0000 00090000 crypt32.dll
76330000 00010000 zcorem.dll
76340000 00010000 winsta.dll
76360000 00010000 msimg32.dll
76370000 00020000 imm32.dll
76390000 00050000 comdlg32.dll
763e0000 00200000 msi.dll
765e0000 00020000 cscdll.dll
76600000 00050000 cscui.dll
76660000 000f0000 setupapi.dll
76750000 00010000 mf3216.dll
76760000 00010000 dnsrslvr.dll
76770000 00010000 shfolder.dll
76780000 00010000 cryptdll.dll
76790000 00020000 ntdsapi.dll
767b0000 00030000 w32time.dll
767e0000 00030000 schannel.dll
76810000 00020000 hlink.dll
76830000 00040000 unidrvui.dll
76870000 00040000 unidrv.dll
768c0000 000b0000 pcl5eres.dll
76970000 00010000 linkinfo.dll
76980000 00030000 ntshrui.dll
769b0000 00150000 shdocvw.dll
76b00000 00010000 ctwdm32.dll
76b10000 00020000 atl.dll
76b30000 00030000 winmm.dll
76b60000 00040000 es.dll
76ba0000 00010000 sfc.dll
76bb0000 00010000 regapi.dll
76bc0000 00020000 shsvcs.dll
76be0000 00010000 psapi.dll
76bf0000 00030000 credui.dll
76c20000 00030000 wintrust.dll
76c50000 00030000 sfc_os.dll
76c80000 00030000 imagehlp.dll
76cb0000 00010000 authz.dll
76cd0000 00020000 ntmarta.dll
76d00000 00020000 msv1_0.dll
76d20000 00010000 wmi.dll
76d30000 00020000 mprapi.dll
76d50000 00020000 iphlpapi.dll
76d70000 00020000 dhcpcsvc.dll
76d90000 00040000 wuaueng.dll
76dd0000 00030000 netman.dll
76e00000 00030000 adsldpc.dll
76e30000 00030000 activeds.dll
76e70000 00010000 rtutils.dll
76e80000 00020000 rasman.dll
76ea0000 00030000 tapi32.dll
76ed0000 00040000 rasapi32.dll
76f10000 00030000 dnsapi.dll
76f40000 00010000 wtsapi32.dll
76f50000 00030000 wldap32.dll
76f80000 00010000 secur32.dll
76fa0000 00010000 winrnr.dll
76fb0000 00010000 rasadhlp.dll
76fc0000 00080000 clbcatq.dll
77040000 000d0000 comres.dll
77110000 00090000 oleaut32.dll
771a0000 00120000 ole32.dll
772c0000 00070000 shlwapi.dll
773c0000 00800000 shell32.dll
77bc0000 00010000 midimap.dll
77bd0000 00020000 msacm32.dll
77bf0000 00010000 version.dll
77c00000 00060000 msvcrt.dll
77c60000 00040000 gdi32.dll
77d30000 00090000 user32.dll
77dc0000 000a0000 advapi32.dll
77e60000 000f0000 kernel32.dll
77f50000 000b0000 ntdll.dll
78000000 00090000 rpcrt4.dll
78190000 001b0000 asms\10100\msft\windows\gdiplus\gdiplus.dll
7c000000 00130000 msvidctl.dll
7c130000 00160000 query.dll
7c290000 001e0000 acgenral.dll
7d650000 00010000 ntvdm64.dll
7d670000 00010000 kbdurs.dll
7d740000 00010000 kbdinori.dll
7d760000 00010000 kbdinmal.dll
7d7b0000 00010000 kbdinben.dll
7d7c0000 00010000 kbdinasa.dll
7d7d0000 00010000 kbdhebx.dll
7d850000 00010000 isetuc0c.dll
7d860000 00010000 isetu816.dll
7d870000 00010000 isetu804.dll
7d880000 00010000 isetu416.dll
7d890000 00010000 isetu40c.dll
7d8a0000 00010000 isetu404.dll
7d8b0000 00010000 isetu02d.dll
7d8c0000 00010000 isetu024.dll
7d8d0000 00010000 isetu021.dll
7d8e0000 00010000 isetu01f.dll
7d8f0000 00010000 isetu01e.dll
7d900000 00010000 isetu01d.dll
7d910000 00010000 isetu01b.dll
7d920000 00010000 isetu01a.dll
7d930000 00010000 isetu019.dll
7d940000 00010000 isetu015.dll
7d950000 00010000 isetu014.dll
7d960000 00010000 isetu013.dll
7d970000 00010000 isetu012.dll
7d980000 00010000 isetu011.dll
7d990000 00010000 isetu010.dll
7d9a0000 00010000 isetu00e.dll
7d9b0000 00010000 isetu00b.dll
7d9c0000 00010000 isetu00a.dll
7d9d0000 00010000 isetu009.dll
7d9e0000 00010000 isetu008.dll
7d9f0000 00010000 isetu007.dll
7da00000 00010000 isetu006.dll
7da10000 00010000 isetu005.dll
7da20000 00010000 isetu003.dll
7da40000 00010000 _setup.dll
7DAE0000 00070000 wow6432\imm32.dll
7DB50000 00060000 wow6432\secur32.dll
7DBB0000 00090000 wow6432\gdi32.dll
7DC40000 000d0000 wow6432\rpcrt4.dll
7DD10000 000d0000 wow6432\user32.dll
7DDE0000 00120000 wow6432\kernel32.dll
7DF00000 00100000 wow6432\ntdll.dll
bfdd0000 001b0000 g400d.dll
bfdd0000 001b0000 nv4.dll
bfed0000 000b0000 3dfxvs.dll
bfee0000 00090000 i81xdnt5.dll
bff00000 00080000 g200d.dll
bff10000 00060000 sgiul50.dll
bff10000 00070000 tridkb.dll
bff20000 00060000 atidrab.dll
bff20000 00060000 atidvag.dll
bff20000 00060000 banshee.dll
bff20000 00060000 i740dnt5.dll
bff30000 00050000 ati2draa.dll
bff30000 00050000 atidvai.dll
bff30000 00050000 trid3d.dll
bff40000 00040000 mgaud.dll
bff40000 00040000 perm2dll.dll
bff40000 00040000 perm3dd.dll
bff40000 00040000 s3mvirge.dll
bff40000 00040000 s3nb.dll
bff40000 00040000 s3sav4.dll
bff40000 00040000 s3savmx.dll
bff40000 00040000 sis300iv.dll
bff50000 00020000 nv3.dll
bff50000 00030000 atidrae.dll
bff50000 00030000 cl546x.dll
bff50000 00030000 s3mt3d.dll
bff50000 00030000 s3sav3d.dll
bff50000 00030000 sis6306v.dll
bff50000 00030000 sisv256.dll
bff50000 00030000 smidispb.dll
bff50000 00030000 t2r4disp.dll
bff60000 00010000 n9i128v2.dll
bff60000 00010000 neo20xx.dll
bff60000 00010000 s3mtrio.dll
bff60000 00020000 ati.dll
bff60000 00020000 atiraged.dll
bff60000 00020000 cirrus.dll
bff60000 00020000 cl5465.dll
bff60000 00020000 n9i3disp.dll
bff60000 00020000 s3legacy.dll
bff60000 00020000 tgiul50.dll
bff70000 00010000 8514a.dll
bff70000 00010000 framebuf.dll
bff70000 00010000 n9i128.dll
bff70000 00010000 vga.dll
bff70000 00010000 vga256.dll
bff70000 00010000 vga64k.dll
bff70000 00010000 w32.dll
bff70000 00010000 weitekp9.dll
bff80000 00020000 dxg.sys
bffa0000 00050000 atmfd.dll
78090000 000f0000 asms\60100\msft\windows\common\controls\comctl32.dll
